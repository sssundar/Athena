magic
tech scmos
timestamp 1434142375
<< polysilicon >>
rect 9 46 35 47
rect 11 45 35 46
rect 7 27 9 39
rect 2 26 9 27
rect -11 23 0 25
rect 4 25 9 26
rect 7 21 14 23
rect 22 21 24 23
rect 7 15 9 21
rect -2 13 0 15
rect 4 13 9 15
rect 11 13 14 15
rect 22 13 24 15
rect 11 11 13 13
rect -2 9 0 11
rect 4 9 13 11
rect -2 5 0 7
rect 4 5 14 7
rect 22 5 24 7
rect -2 -3 0 -1
rect 4 -3 14 -1
rect 22 -3 24 -1
rect -2 -7 0 -5
rect 4 -7 13 -5
rect 11 -9 13 -7
rect -2 -11 0 -9
rect 4 -11 9 -9
rect 11 -11 14 -9
rect 22 -11 24 -9
rect 7 -17 9 -11
rect -18 -21 0 -19
rect 7 -19 14 -17
rect 22 -19 24 -17
rect 2 -25 4 -22
rect 2 -27 8 -25
rect 6 -35 8 -27
rect 11 -42 41 -41
rect 9 -43 41 -42
<< ndiffusion >>
rect 0 15 4 16
rect 0 11 4 13
rect 0 7 4 9
rect 0 4 4 5
rect 0 -1 4 0
rect 0 -5 4 -3
rect 0 -9 4 -7
rect 0 -12 4 -11
<< pdiffusion >>
rect 14 23 22 24
rect 14 20 22 21
rect 14 15 22 16
rect 14 12 22 13
rect 14 7 22 8
rect 14 4 22 5
rect 14 -1 22 0
rect 14 -4 22 -3
rect 14 -9 22 -8
rect 14 -12 22 -11
rect 14 -17 22 -16
rect 14 -20 22 -19
<< metal1 >>
rect -7 36 -4 47
rect 29 36 32 47
rect -7 32 0 36
rect 22 32 32 36
rect -22 -43 -19 -22
rect -15 -43 -12 22
rect -7 -43 -4 32
rect 0 20 4 22
rect 7 24 14 27
rect 7 20 10 24
rect 29 20 32 32
rect 4 17 10 20
rect 7 12 10 17
rect 22 16 32 20
rect 7 9 14 12
rect 29 4 32 16
rect 22 0 32 4
rect 7 -8 14 -5
rect 7 -13 10 -8
rect 29 -12 32 0
rect 4 -16 10 -13
rect 22 -16 32 -12
rect 0 -18 4 -16
rect 7 -20 10 -16
rect 7 -23 14 -20
rect 29 -43 32 -16
rect 35 -43 38 43
<< ntransistor >>
rect 0 13 4 15
rect 0 9 4 11
rect 0 5 4 7
rect 0 -3 4 -1
rect 0 -7 4 -5
rect 0 -11 4 -9
<< ptransistor >>
rect 14 21 22 23
rect 14 13 22 15
rect 14 5 22 7
rect 14 -3 22 -1
rect 14 -11 22 -9
rect 14 -19 22 -17
<< polycontact >>
rect 7 42 11 46
rect 35 43 39 47
rect -15 22 -11 26
rect 0 22 4 26
rect -22 -22 -18 -18
rect 0 -22 4 -18
rect 7 -42 11 -38
rect 41 -43 45 -39
<< ndcontact >>
rect 0 16 4 20
rect 0 0 4 4
rect 0 -16 4 -12
<< pdcontact >>
rect 14 24 22 28
rect 14 16 22 20
rect 14 8 22 12
rect 14 0 22 4
rect 14 -8 22 -4
rect 14 -16 22 -12
rect 14 -24 22 -20
use inverter  inverter_0
timestamp 1430424850
transform 0 1 -7 1 0 37
box -5 5 7 31
use inverter  inverter_1
timestamp 1430424850
transform 0 1 -7 -1 0 -33
box -5 5 7 31
<< labels >>
rlabel metal1 -22 -24 -19 -22 3 w
rlabel metal1 35 -24 38 -22 1 r_
rlabel metal1 -7 -24 -4 -22 1 GND
rlabel metal1 29 -24 32 -22 1 Vdd
rlabel metal1 -15 -24 -12 -22 1 r
rlabel polycontact 42 -43 45 -40 8 w_
rlabel polysilicon 23 -18 23 -18 1 regw
rlabel polysilicon 23 -10 23 -10 1 phi0
rlabel polysilicon 23 -2 23 -2 1 wr_id
rlabel polysilicon 23 6 23 6 1 rd_id
rlabel polysilicon 23 14 23 14 1 phi1
rlabel polysilicon 23 22 23 22 1 regr
<< end >>
