magic
tech scmos
timestamp 1434158754
<< polysilicon >>
rect -16 37 -14 49
rect -8 37 -6 52
rect 8 37 10 52
rect 16 37 18 52
rect 32 37 34 52
rect -24 33 -23 37
rect -25 31 -23 33
rect -25 29 -19 31
rect -21 14 -19 29
rect -16 25 -14 33
rect -8 29 -6 33
rect -8 27 3 29
rect -16 23 -1 25
rect -3 21 -1 23
rect 1 21 3 27
rect 8 25 10 33
rect 16 30 18 33
rect 16 28 26 30
rect 8 23 22 25
rect 20 21 22 23
rect 24 21 26 28
rect 32 21 34 33
rect -21 12 -16 14
rect -32 -2 -30 12
rect -34 -4 -28 -2
rect -20 -4 -18 -2
rect -34 -10 -32 -4
rect -16 -6 -14 12
rect -3 9 -1 11
rect 1 9 3 11
rect 20 9 22 11
rect 24 9 26 11
rect 32 9 34 11
rect -30 -8 -28 -6
rect -20 -8 -14 -6
rect -12 0 -8 2
rect -12 -7 -10 0
rect -34 -12 -29 -10
rect -31 -28 -29 -12
rect -19 -14 -17 -8
rect -23 -16 -17 -14
rect -12 -9 -8 -7
rect -23 -23 -21 -16
rect -12 -18 -10 -9
rect 40 0 44 2
rect 42 -7 44 0
rect 40 -9 44 -7
rect -12 -20 -7 -18
rect -3 -20 9 -18
rect 18 -18 25 -16
rect 42 -18 44 -9
rect 7 -22 9 -20
rect 23 -20 44 -18
rect 23 -22 25 -20
rect -31 -30 -25 -28
rect -23 -29 -21 -27
rect -27 -31 -25 -30
rect -27 -37 -25 -35
rect 7 -40 9 -38
rect 23 -40 25 -38
<< ndiffusion >>
rect -17 33 -16 37
rect -14 33 -13 37
rect -9 33 -8 37
rect -6 33 -5 37
rect 7 33 8 37
rect 10 33 11 37
rect 15 33 16 37
rect 18 33 19 37
rect 31 33 32 37
rect 34 33 35 37
rect -24 -27 -23 -23
rect -21 -27 -20 -23
rect -28 -35 -27 -31
rect -25 -35 -24 -31
rect 6 -38 7 -22
rect 9 -38 10 -22
rect 22 -38 23 -22
rect 25 -38 26 -22
<< pdiffusion >>
rect -28 -2 -20 -1
rect -28 -6 -20 -4
rect -4 11 -3 21
rect -1 11 1 21
rect 3 11 4 21
rect 19 11 20 21
rect 22 11 24 21
rect 26 11 27 21
rect 31 11 32 21
rect 34 11 35 21
rect -8 2 10 5
rect -8 -1 7 0
rect 6 -6 7 -1
rect -8 -7 7 -6
rect -28 -9 -20 -8
rect 9 -9 10 2
rect -8 -12 10 -9
rect 22 2 40 5
rect 22 -9 23 2
rect 25 -1 40 0
rect 25 -6 26 -1
rect 25 -7 40 -6
rect 22 -12 40 -9
<< metal1 >>
rect -4 46 39 49
rect -4 44 -1 46
rect -21 41 -1 44
rect -21 37 -18 41
rect -4 37 -1 41
rect -24 33 -21 37
rect 3 40 23 43
rect 3 37 6 40
rect 20 37 23 40
rect 35 37 39 46
rect 23 33 27 37
rect -12 30 -9 33
rect 10 30 15 33
rect -35 27 13 30
rect 7 26 12 27
rect 16 24 39 27
rect 15 21 19 24
rect 36 21 39 24
rect -12 12 -8 16
rect 8 11 15 21
rect 27 8 31 11
rect -34 5 44 8
rect -28 3 -20 5
rect -28 -17 -24 -13
rect 2 -15 6 -6
rect -28 -20 -7 -17
rect 2 -19 14 -15
rect -28 -23 -24 -20
rect 2 -22 6 -19
rect 26 -22 30 -6
rect -31 -31 -28 -23
rect -20 -40 -17 -27
rect -34 -44 -20 -41
rect 2 -47 6 -38
rect 14 -40 18 -38
rect 26 -47 30 -38
rect 41 -44 44 -41
<< metal2 >>
rect -16 -44 14 -41
rect 18 -44 37 -41
<< ntransistor >>
rect -16 33 -14 37
rect -8 33 -6 37
rect 8 33 10 37
rect 16 33 18 37
rect 32 33 34 37
rect -23 -27 -21 -23
rect -27 -35 -25 -31
rect 7 -38 9 -22
rect 23 -38 25 -22
<< ptransistor >>
rect -28 -4 -20 -2
rect -3 11 -1 21
rect 1 11 3 21
rect 20 11 22 21
rect 24 11 26 21
rect 32 11 34 21
rect -28 -8 -20 -6
rect -8 0 9 2
rect 7 -7 9 0
rect -8 -9 9 -7
rect 23 0 40 2
rect 23 -7 25 0
rect 23 -9 40 -7
<< polycontact >>
rect -18 49 -14 53
rect -8 52 -4 56
rect 6 52 10 56
rect 16 52 20 56
rect 30 52 34 56
rect -28 33 -24 37
rect -32 12 -28 16
rect -16 12 -12 16
rect -7 -20 -3 -16
rect 14 -19 18 -15
<< ndcontact >>
rect -21 33 -17 37
rect -13 33 -9 37
rect -5 33 -1 37
rect 3 33 7 37
rect 11 33 15 37
rect 19 33 23 37
rect 27 33 31 37
rect 35 33 39 37
rect -28 -27 -24 -23
rect -20 -27 -16 -23
rect -32 -35 -28 -31
rect -24 -35 -20 -31
rect 2 -38 6 -22
rect 10 -38 14 -22
rect 18 -38 22 -22
rect 26 -38 30 -22
<< pdcontact >>
rect -28 -1 -20 3
rect -8 11 -4 21
rect 4 11 8 21
rect 15 11 19 21
rect 27 11 31 21
rect 35 11 39 21
rect -8 -6 6 -1
rect -28 -13 -20 -9
rect 10 -12 14 5
rect 18 -12 22 5
rect 26 -6 40 -1
<< m2contact >>
rect -20 -44 -16 -40
rect 14 -44 18 -40
rect 37 -44 41 -40
<< psubstratepcontact >>
rect 14 -38 18 -22
<< nsubstratencontact >>
rect 14 -12 18 5
<< labels >>
rlabel metal1 -11 6 -11 6 5 Vdd
rlabel polycontact 14 -16 14 -16 1 read_
rlabel metal1 28 -16 28 -16 1 read
rlabel polycontact -16 15 -16 15 5 ungatedRead_
rlabel metal1 -33 29 -33 29 3 GND
rlabel polycontact -32 16 -32 16 4 phi1_
rlabel polycontact -16 51 -16 51 5 instructionCycleCountIs0
rlabel polycontact -6 54 -6 54 5 instructionCycleCountIs2
rlabel polycontact 8 54 8 54 5 BranchInstruction
rlabel polycontact 18 54 18 54 5 InputInstruction
rlabel polycontact 32 54 32 54 5 instructionCycleCountIs1
<< end >>
