magic
tech scmos
timestamp 1433954011
<< polysilicon >>
rect 58 68 60 70
rect 28 24 32 26
rect 28 -18 30 24
rect 66 1 104 3
rect 74 -5 104 -3
rect 42 -8 48 -6
rect 56 -8 59 -6
rect 42 -10 44 -8
rect 32 -12 34 -10
rect 38 -12 44 -10
rect 57 -10 64 -8
rect 42 -16 48 -14
rect 56 -16 58 -14
rect 42 -18 44 -16
rect 28 -20 34 -18
rect 38 -20 44 -18
rect 62 -17 64 -10
rect 32 -24 34 -22
rect 38 -24 48 -22
rect 56 -24 59 -22
rect 74 -24 76 -5
rect 57 -26 76 -24
<< ndiffusion >>
rect 34 -10 38 -9
rect 34 -13 38 -12
rect 34 -18 38 -17
rect 34 -22 38 -20
rect 34 -25 38 -24
<< pdiffusion >>
rect 48 -6 56 -5
rect 48 -9 56 -8
rect 48 -14 56 -13
rect 48 -17 56 -16
rect 48 -22 56 -21
rect 48 -25 56 -24
<< metal1 >>
rect 0 85 3 88
rect 7 85 10 88
rect 14 85 17 88
rect 21 85 24 88
rect 28 85 31 88
rect 70 85 73 88
rect 77 85 80 88
rect 84 85 87 88
rect 91 85 94 88
rect 98 85 101 88
rect 41 35 45 38
rect 105 5 108 88
rect 0 -29 3 0
rect 7 -29 10 0
rect 14 -29 17 0
rect 21 -29 24 0
rect 28 -13 31 0
rect 41 -5 48 -2
rect 56 -4 66 -1
rect 38 -8 44 -5
rect 70 -9 73 0
rect 56 -13 73 -9
rect 28 -17 34 -13
rect 28 -29 31 -17
rect 41 -21 48 -17
rect 56 -21 62 -17
rect 41 -25 45 -21
rect 70 -25 73 -13
rect 38 -29 45 -25
rect 56 -29 73 -25
rect 77 -29 80 0
rect 84 -29 87 0
rect 91 -29 94 0
rect 98 -29 101 0
rect 105 -29 108 -7
<< ntransistor >>
rect 34 -12 38 -10
rect 34 -20 38 -18
rect 34 -24 38 -22
<< ptransistor >>
rect 48 -8 56 -6
rect 48 -16 56 -14
rect 48 -24 56 -22
<< polycontact >>
rect 62 -1 66 3
rect 104 1 108 5
rect 62 -21 66 -17
rect 104 -7 108 -3
<< ndcontact >>
rect 34 -9 38 -5
rect 34 -17 38 -13
rect 34 -29 38 -25
<< pdcontact >>
rect 48 -5 56 -1
rect 48 -13 56 -9
rect 48 -21 56 -17
rect 48 -29 56 -25
<< m2contact >>
rect 41 84 45 88
use accumbit  accumbit_0
timestamp 1433920747
transform 1 0 35 0 1 69
box -35 -69 66 19
<< labels >>
rlabel metal1 105 -29 108 -26 8 zin
rlabel metal1 105 85 108 88 6 zout
rlabel metal1 0 85 3 88 4 phi1
rlabel metal1 7 85 10 88 5 ld
rlabel metal1 14 85 17 88 5 w
rlabel metal1 21 85 24 88 5 r
rlabel m2contact 41 84 45 88 5 bus
rlabel metal1 28 85 31 88 5 GND
rlabel metal1 70 85 73 88 5 Vdd
rlabel metal1 77 85 80 88 5 r_
rlabel metal1 84 85 87 88 5 w_
rlabel metal1 91 85 94 88 5 ld_
rlabel metal1 98 85 101 88 5 phi1_
rlabel polysilicon 59 69 59 69 1 in
rlabel metal1 41 35 45 38 1 out
<< end >>
