magic
tech scmos
timestamp 1434158463
<< polysilicon >>
rect 23 17 25 19
rect -15 5 -1 7
rect 25 5 44 7
rect -8 -3 -1 -1
rect 25 -3 37 -1
rect -29 -15 1 -13
rect 5 -15 7 -13
rect 12 -15 14 -5
rect 12 -17 19 -15
rect -22 -35 -1 -33
rect 9 -44 11 -31
rect 25 -35 51 -33
rect 9 -46 26 -44
rect 24 -56 26 -46
<< ndiffusion >>
rect 1 -13 5 -12
rect 1 -16 5 -15
<< metal1 >>
rect -33 -12 -30 24
rect -33 -75 -30 -16
rect -26 -32 -23 24
rect -19 8 -16 24
rect -26 -75 -23 -36
rect -19 -75 -16 4
rect -12 0 -9 24
rect -5 16 -2 24
rect -5 12 1 16
rect 8 14 12 20
rect 31 16 34 24
rect -12 -75 -9 -4
rect -5 -8 -2 12
rect 23 12 34 16
rect -5 -12 1 -8
rect -5 -24 -2 -12
rect 8 -16 11 2
rect 31 -8 34 12
rect 38 0 41 24
rect 45 8 48 24
rect 23 -12 34 -8
rect 5 -20 11 -16
rect -5 -28 1 -24
rect 8 -25 11 -20
rect 31 -24 34 -12
rect -5 -63 -2 -28
rect 23 -28 34 -24
rect 11 -40 15 -37
rect 31 -63 34 -28
rect -5 -67 1 -63
rect 29 -67 34 -63
rect -5 -75 -2 -67
rect 31 -75 34 -67
rect 38 -75 41 -4
rect 45 -75 48 4
rect 52 -32 55 24
rect 52 -75 55 -36
<< ntransistor >>
rect 1 -15 5 -13
<< polycontact >>
rect 8 10 12 14
rect -19 4 -15 8
rect 44 4 48 8
rect -12 -4 -8 0
rect 37 -4 41 0
rect -33 -16 -29 -12
rect 19 -19 23 -15
rect 8 -29 12 -25
rect -26 -36 -22 -32
rect 51 -36 55 -32
<< ndcontact >>
rect 1 -12 5 -8
rect 1 -20 5 -16
use inverter  inverter_0
timestamp 1430424850
transform 0 1 -6 1 0 17
box -5 5 7 31
use latch  latch_0
timestamp 1430426212
transform 0 1 1 -1 0 10
box -6 -2 10 24
use latch  latch_1
timestamp 1430426212
transform 0 1 1 1 0 -6
box -6 -2 10 24
use latch  latch_2
timestamp 1430426212
transform 0 1 1 -1 0 -30
box -6 -2 10 24
use staticizer  staticizer_0
timestamp 1430428783
transform 0 1 -3 -1 0 -63
box -19 2 12 32
<< labels >>
rlabel polycontact 21 -17 21 -17 8 inc_in
rlabel metal1 11 -40 14 -37 1 inc_out
rlabel metal1 8 -20 11 -17 1 addr_out
rlabel metal1 -5 21 -2 24 5 GND
rlabel metal1 31 21 34 24 6 Vdd
rlabel polysilicon 24 18 24 18 1 branch_in
rlabel metal1 -12 21 -9 24 4 inc_w
rlabel metal1 38 21 41 24 5 inc_w_
rlabel metal1 45 21 48 24 5 branch_w_
rlabel metal1 -19 21 -16 24 5 branch_w
rlabel metal1 -26 21 -23 24 5 phi1
rlabel metal1 52 21 55 24 6 phi1_
rlabel metal1 -33 21 -30 24 4 reset
<< end >>
