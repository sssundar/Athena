magic
tech scmos
timestamp 1434090485
<< polysilicon >>
rect -67 -111 -65 -102
rect -59 -111 -57 -102
rect -17 -111 -15 -102
rect -9 -111 -7 -102
rect 7 -111 9 -102
rect 33 -111 35 -102
rect 41 -111 43 -102
rect 57 -111 59 -102
rect -89 -125 -75 -123
rect -89 -146 -87 -125
rect -67 -125 -65 -119
rect -59 -125 -57 -119
rect -67 -127 -63 -125
rect -65 -129 -63 -127
rect -61 -127 -57 -125
rect -31 -125 -24 -123
rect -61 -129 -59 -127
rect -65 -135 -63 -133
rect -61 -135 -59 -133
rect -89 -148 -85 -146
rect -89 -155 -87 -148
rect -89 -157 -85 -155
rect -89 -166 -87 -157
rect -31 -146 -29 -125
rect -17 -125 -15 -119
rect -9 -121 -7 -119
rect -9 -123 -2 -121
rect -17 -127 -6 -125
rect -8 -129 -6 -127
rect -4 -129 -2 -123
rect 7 -125 9 -119
rect 0 -127 9 -125
rect 0 -129 2 -127
rect -8 -135 -6 -133
rect -4 -135 -2 -133
rect 0 -135 2 -133
rect -37 -148 -33 -146
rect -35 -155 -33 -148
rect -37 -157 -33 -155
rect -89 -168 -68 -166
rect -59 -166 -52 -164
rect -35 -166 -33 -157
rect -70 -170 -68 -168
rect -54 -168 -33 -166
rect -31 -148 -27 -146
rect -31 -155 -29 -148
rect -31 -157 -27 -155
rect -31 -166 -29 -157
rect 27 -146 29 -126
rect 33 -125 35 -119
rect 41 -121 43 -119
rect 41 -123 48 -121
rect 33 -127 44 -125
rect 42 -129 44 -127
rect 46 -129 48 -123
rect 57 -125 59 -119
rect 50 -127 59 -125
rect 50 -129 52 -127
rect 42 -135 44 -133
rect 46 -135 48 -133
rect 50 -135 52 -133
rect 21 -148 25 -146
rect 23 -155 25 -148
rect 21 -157 25 -155
rect -31 -168 -10 -166
rect -1 -166 6 -164
rect 23 -166 25 -157
rect -54 -170 -52 -168
rect -12 -170 -10 -168
rect 4 -168 25 -166
rect 27 -148 31 -146
rect 27 -155 29 -148
rect 27 -157 31 -155
rect 27 -166 29 -157
rect 79 -148 83 -146
rect 81 -155 83 -148
rect 79 -157 83 -155
rect 27 -168 48 -166
rect 57 -166 64 -164
rect 81 -166 83 -157
rect 4 -170 6 -168
rect 46 -170 48 -168
rect 62 -168 83 -166
rect 62 -170 64 -168
rect -70 -188 -68 -186
rect -54 -188 -52 -186
rect -12 -188 -10 -186
rect 4 -188 6 -186
rect 46 -188 48 -186
rect 62 -188 64 -186
<< ndiffusion >>
rect -66 -133 -65 -129
rect -63 -133 -61 -129
rect -59 -133 -58 -129
rect -9 -133 -8 -129
rect -6 -133 -4 -129
rect -2 -133 0 -129
rect 2 -133 3 -129
rect 41 -133 42 -129
rect 44 -133 46 -129
rect 48 -133 50 -129
rect 52 -133 53 -129
rect -71 -186 -70 -170
rect -68 -186 -67 -170
rect -55 -186 -54 -170
rect -52 -186 -51 -170
rect -13 -186 -12 -170
rect -10 -186 -9 -170
rect 3 -186 4 -170
rect 6 -186 7 -170
rect 45 -186 46 -170
rect 48 -186 49 -170
rect 61 -186 62 -170
rect 64 -186 65 -170
<< pdiffusion >>
rect -68 -119 -67 -111
rect -65 -119 -64 -111
rect -60 -119 -59 -111
rect -57 -119 -56 -111
rect -18 -119 -17 -111
rect -15 -119 -14 -111
rect -10 -119 -9 -111
rect -7 -119 -6 -111
rect 6 -119 7 -111
rect 9 -119 10 -111
rect 32 -119 33 -111
rect 35 -119 36 -111
rect 40 -119 41 -111
rect 43 -119 44 -111
rect 56 -119 57 -111
rect 59 -119 60 -111
rect -85 -146 -67 -143
rect -85 -149 -70 -148
rect -71 -154 -70 -149
rect -85 -155 -70 -154
rect -68 -157 -67 -146
rect -85 -160 -67 -157
rect -55 -146 -37 -143
rect -27 -146 -9 -143
rect -55 -157 -54 -146
rect -52 -149 -37 -148
rect -52 -154 -51 -149
rect -52 -155 -37 -154
rect -55 -160 -37 -157
rect -27 -149 -12 -148
rect -13 -154 -12 -149
rect -27 -155 -12 -154
rect -10 -157 -9 -146
rect -27 -160 -9 -157
rect 3 -146 21 -143
rect 31 -146 49 -143
rect 3 -157 4 -146
rect 6 -149 21 -148
rect 6 -154 7 -149
rect 6 -155 21 -154
rect 3 -160 21 -157
rect 31 -149 46 -148
rect 45 -154 46 -149
rect 31 -155 46 -154
rect 48 -157 49 -146
rect 31 -160 49 -157
rect 61 -146 79 -143
rect 61 -157 62 -146
rect 64 -149 79 -148
rect 64 -154 65 -149
rect 64 -155 79 -154
rect 61 -160 79 -157
<< metal1 >>
rect -55 -102 -17 -98
rect -89 -108 83 -105
rect -64 -111 -61 -108
rect -14 -111 -10 -108
rect 10 -111 18 -108
rect 36 -111 40 -108
rect 60 -111 64 -108
rect -72 -122 -69 -119
rect -55 -122 -52 -119
rect -22 -122 -19 -119
rect -5 -122 -2 -119
rect 2 -122 5 -119
rect 28 -122 31 -119
rect 45 -122 48 -119
rect 52 -122 55 -119
rect -71 -125 -52 -122
rect -71 -126 -69 -125
rect -20 -125 5 -122
rect -72 -129 -69 -126
rect -13 -129 -9 -125
rect 29 -125 55 -122
rect 37 -129 41 -125
rect -91 -133 -79 -129
rect -72 -133 -70 -129
rect -54 -133 -53 -129
rect 11 -133 12 -129
rect 57 -133 58 -129
rect -91 -188 -88 -133
rect 80 -140 83 -108
rect -85 -143 83 -140
rect -75 -163 -71 -154
rect -75 -167 -63 -163
rect -75 -170 -71 -167
rect -51 -170 -47 -154
rect -17 -163 -13 -154
rect -17 -167 -5 -163
rect -17 -170 -13 -167
rect 7 -170 11 -154
rect 41 -163 45 -154
rect 41 -167 53 -163
rect 41 -170 45 -167
rect 65 -170 69 -154
rect -63 -188 -59 -186
rect -5 -188 -1 -186
rect 53 -188 57 -186
rect 76 -192 83 -189
<< metal2 >>
rect -75 -133 -53 -129
rect -49 -133 7 -129
rect 16 -133 58 -129
rect -87 -192 -63 -189
rect -59 -192 -5 -189
rect -1 -192 53 -189
rect 57 -192 72 -189
<< ntransistor >>
rect -65 -133 -63 -129
rect -61 -133 -59 -129
rect -8 -133 -6 -129
rect -4 -133 -2 -129
rect 0 -133 2 -129
rect 42 -133 44 -129
rect 46 -133 48 -129
rect 50 -133 52 -129
rect -70 -186 -68 -170
rect -54 -186 -52 -170
rect -12 -186 -10 -170
rect 4 -186 6 -170
rect 46 -186 48 -170
rect 62 -186 64 -170
<< ptransistor >>
rect -67 -119 -65 -111
rect -59 -119 -57 -111
rect -17 -119 -15 -111
rect -9 -119 -7 -111
rect 7 -119 9 -111
rect 33 -119 35 -111
rect 41 -119 43 -111
rect 57 -119 59 -111
rect -85 -148 -68 -146
rect -70 -155 -68 -148
rect -85 -157 -68 -155
rect -54 -148 -37 -146
rect -54 -155 -52 -148
rect -54 -157 -37 -155
rect -27 -148 -10 -146
rect -12 -155 -10 -148
rect -27 -157 -10 -155
rect 4 -148 21 -146
rect 4 -155 6 -148
rect 4 -157 21 -155
rect 31 -148 48 -146
rect 46 -155 48 -148
rect 31 -157 48 -155
rect 62 -148 79 -146
rect 62 -155 64 -148
rect 62 -157 79 -155
<< polycontact >>
rect -69 -102 -65 -98
rect -59 -102 -55 -98
rect -17 -102 -13 -98
rect -9 -102 -5 -98
rect 5 -102 9 -98
rect 33 -102 37 -98
rect 41 -102 45 -98
rect 55 -102 59 -98
rect -75 -126 -71 -122
rect -24 -126 -20 -122
rect 25 -126 29 -122
rect -63 -167 -59 -163
rect -5 -167 -1 -163
rect 53 -167 57 -163
<< ndcontact >>
rect -70 -133 -66 -129
rect -58 -133 -54 -129
rect -13 -133 -9 -129
rect 3 -133 7 -129
rect 37 -133 41 -129
rect 53 -133 57 -129
rect -75 -186 -71 -170
rect -67 -186 -63 -170
rect -59 -186 -55 -170
rect -51 -186 -47 -170
rect -17 -186 -13 -170
rect -9 -186 -5 -170
rect -1 -186 3 -170
rect 7 -186 11 -170
rect 41 -186 45 -170
rect 49 -186 53 -170
rect 57 -186 61 -170
rect 65 -186 69 -170
<< pdcontact >>
rect -72 -119 -68 -111
rect -64 -119 -60 -111
rect -56 -119 -52 -111
rect -22 -119 -18 -111
rect -14 -119 -10 -111
rect -6 -119 -2 -111
rect 2 -119 6 -111
rect 10 -119 14 -111
rect 28 -119 32 -111
rect 36 -119 40 -111
rect 44 -119 48 -111
rect 52 -119 56 -111
rect 60 -119 64 -111
rect -85 -154 -71 -149
rect -67 -160 -63 -143
rect -59 -160 -55 -143
rect -51 -154 -37 -149
rect -27 -154 -13 -149
rect -9 -160 -5 -143
rect -1 -160 3 -143
rect 7 -154 21 -149
rect 31 -154 45 -149
rect 49 -160 53 -143
rect 57 -160 61 -143
rect 65 -154 79 -149
<< m2contact >>
rect -79 -133 -75 -129
rect -53 -133 -49 -129
rect 12 -133 16 -129
rect 58 -133 62 -129
rect -91 -192 -87 -188
rect -63 -192 -59 -188
rect -5 -192 -1 -188
rect 53 -192 57 -188
rect 72 -192 76 -188
<< psubstratepcontact >>
rect 7 -133 11 -129
rect -63 -186 -59 -170
rect -5 -186 -1 -170
rect 53 -186 57 -170
<< nsubstratencontact >>
rect 14 -119 18 -111
rect -63 -160 -59 -143
rect -5 -160 -1 -143
rect 53 -160 57 -143
<< labels >>
rlabel metal1 -38 -100 -38 -100 5 phi0
rlabel polycontact -67 -100 -67 -100 5 ArithmeticInstruction
rlabel polycontact -7 -100 -7 -100 5 simpleWrite
rlabel polycontact 7 -100 7 -100 5 Register0Write
rlabel polycontact 35 -100 35 -100 5 phi1
rlabel polycontact 43 -100 43 -100 5 simpleRead
rlabel polycontact 57 -100 57 -100 5 Register0Read
rlabel metal2 -34 -191 -34 -191 1 GND
rlabel metal1 -37 -107 -37 -107 1 Vdd
rlabel metal1 -73 -163 -73 -163 1 writeFromAdder
rlabel metal1 -50 -163 -50 -163 1 writeFromAdder_
rlabel metal1 -15 -164 -15 -164 1 writeFromDP
rlabel metal1 9 -164 9 -164 1 writeFromDP_
rlabel metal1 43 -164 43 -164 1 readToDP
rlabel metal1 67 -164 67 -164 1 readToDP_
<< end >>
