magic
tech scmos
timestamp 1430441829
<< polysilicon >>
rect -2 155 0 157
rect 6 155 8 162
rect -2 120 0 123
rect -1 116 0 120
rect -2 113 0 116
rect 6 113 8 123
rect 15 117 24 119
rect -2 95 0 97
rect 6 95 8 97
rect -9 80 -7 82
rect -3 80 7 82
rect 15 80 17 82
rect -21 71 4 73
rect -2 57 0 59
rect 6 57 8 64
rect -2 22 0 25
rect -1 18 0 22
rect -2 15 0 18
rect 6 15 8 25
rect 15 19 24 21
rect -2 -3 0 -1
rect 6 -3 8 -1
rect -23 -27 4 -25
<< ndiffusion >>
rect -3 97 -2 113
rect 0 97 6 113
rect 8 97 9 113
rect -7 82 -3 83
rect -7 79 -3 80
rect -3 -1 -2 15
rect 0 -1 6 15
rect 8 -1 9 15
<< pdiffusion >>
rect -3 123 -2 155
rect 0 127 6 155
rect 0 123 1 127
rect 5 123 6 127
rect 8 123 9 155
rect 7 82 15 83
rect 7 79 15 80
rect -3 25 -2 57
rect 0 29 6 57
rect 0 25 1 29
rect 5 25 6 29
rect 8 25 9 57
<< metal1 >>
rect -18 93 -15 166
rect 3 162 4 166
rect 18 159 21 166
rect -7 156 21 159
rect -7 155 -3 156
rect 9 155 21 156
rect 17 151 21 155
rect -6 116 -5 120
rect 2 118 5 123
rect 9 118 11 119
rect 2 116 11 118
rect 2 115 12 116
rect 9 113 12 115
rect -5 93 -4 97
rect 9 93 12 97
rect -18 89 -4 93
rect -24 -17 -21 71
rect -33 -20 -21 -17
rect -18 -5 -15 89
rect -7 87 -4 89
rect 1 90 12 93
rect 1 86 4 90
rect 18 89 21 151
rect 19 85 21 89
rect 15 84 21 85
rect -3 77 7 79
rect -3 75 0 77
rect 4 75 7 77
rect 3 64 4 68
rect 18 61 21 84
rect -7 58 21 61
rect -7 57 -3 58
rect 9 57 21 58
rect 17 53 21 57
rect -6 18 -5 22
rect 2 20 5 25
rect 9 20 11 21
rect 2 18 11 20
rect 2 17 12 18
rect 9 15 12 17
rect -5 -5 -4 -1
rect 9 -5 12 -1
rect -18 -9 -4 -5
rect -33 -28 -30 -20
rect -26 -28 -23 -27
rect -18 -28 -15 -9
rect -7 -11 -4 -9
rect 1 -8 12 -5
rect 1 -12 4 -8
rect 18 -9 21 53
rect 24 28 27 116
rect 24 25 34 28
rect 19 -13 21 -9
rect 15 -14 21 -13
rect 18 -28 21 -14
rect 24 -28 27 18
rect 31 -28 34 25
<< ntransistor >>
rect -2 97 0 113
rect 6 97 8 113
rect -7 80 -3 82
rect -2 -1 0 15
rect 6 -1 8 15
<< ptransistor >>
rect -2 123 0 155
rect 6 123 8 155
rect 7 80 15 82
rect -2 25 0 57
rect 6 25 8 57
<< polycontact >>
rect 4 162 8 166
rect -5 116 -1 120
rect 11 116 15 120
rect 24 116 28 120
rect 0 82 4 86
rect -25 71 -21 75
rect 0 73 4 77
rect 4 64 8 68
rect -5 18 -1 22
rect 11 18 15 22
rect 24 18 28 22
rect 0 -16 4 -12
rect -27 -27 -23 -23
rect 0 -25 4 -21
<< ndcontact >>
rect -7 97 -3 113
rect 9 97 13 113
rect -7 83 -3 87
rect -7 75 -3 79
rect -7 -1 -3 15
rect 9 -1 13 15
<< pdcontact >>
rect -7 123 -3 155
rect 1 123 5 127
rect 9 123 13 155
rect 7 83 15 87
rect 7 75 15 79
rect -7 25 -3 57
rect 1 25 5 29
rect 9 25 13 57
<< m2contact >>
rect -1 162 3 166
rect -10 116 -6 120
rect -1 64 3 68
rect -10 18 -6 22
<< psubstratepcontact >>
rect -9 93 -5 97
rect -9 -5 -5 -1
<< nsubstratencontact >>
rect 13 151 17 155
rect 15 85 19 89
rect 13 53 17 57
rect 15 -13 19 -9
use inverter  inverter_0
timestamp 1430424850
transform 0 1 -14 -1 0 -16
box -5 5 7 31
<< labels >>
rlabel metal1 2 77 2 77 1 out
rlabel metal1 -18 -28 -15 -25 1 GND
rlabel metal1 18 -28 21 -25 1 Vdd
rlabel metal1 24 -28 27 -25 1 r_
rlabel metal1 31 -28 34 -25 8 w_
rlabel metal1 -26 -28 -23 -25 1 r
rlabel metal1 -33 -28 -30 -25 2 w
rlabel m2contact -10 18 -6 22 1 phi1
rlabel m2contact -10 116 -6 120 1 phi0
rlabel m2contact -1 64 3 68 1 regr
rlabel m2contact -1 162 3 166 5 regw
<< end >>
