magic
tech scmos
timestamp 1434174658
<< polysilicon >>
rect -15 30 -5 32
rect 27 30 93 32
rect -15 14 -13 30
rect -8 26 -5 28
rect 27 26 29 28
rect -8 20 -6 26
rect -8 18 8 20
rect -15 12 -8 14
rect -10 3 -8 12
rect 6 3 8 18
rect -10 -31 -8 -29
rect 6 -33 8 -29
<< ndiffusion >>
rect -5 32 27 33
rect -5 28 27 30
rect -5 25 27 26
<< pdiffusion >>
rect -11 -29 -10 3
rect -8 -29 -7 3
rect 5 -29 6 3
rect 8 -29 9 3
<< metal1 >>
rect -15 44 49 47
rect -15 17 -12 44
rect 27 37 37 41
rect 34 31 37 37
rect 93 22 97 29
rect -3 17 1 21
rect -15 14 21 17
rect -15 3 -12 14
rect 10 3 13 14
rect 10 -37 95 -34
<< ntransistor >>
rect -5 30 27 32
rect -5 26 27 28
<< ptransistor >>
rect -10 -29 -8 3
rect 6 -29 8 3
<< polycontact >>
rect 93 29 97 33
rect 6 -37 10 -33
<< ndcontact >>
rect -5 33 27 37
rect -5 21 27 25
<< pdcontact >>
rect -15 -29 -11 3
rect -7 -29 -3 3
rect 1 -29 5 3
rect 9 -29 13 3
<< psubstratepcontact >>
rect -5 37 27 41
<< nsubstratencontact >>
rect -3 -29 1 3
<< labels >>
rlabel metal1 20 16 20 16 7 cout
rlabel metal1 47 46 47 46 5 Cin2
<< end >>
