magic
tech scmos
timestamp 1434088956
<< polysilicon >>
rect 0 9 2 11
rect 6 10 9 11
rect 13 10 16 11
rect 6 9 16 10
rect 24 9 26 11
rect 10 -6 12 0
rect -7 -11 0 -9
rect 26 -11 33 -9
<< ndiffusion >>
rect 2 11 6 12
rect 2 8 6 9
<< pdiffusion >>
rect 16 11 24 12
rect 16 8 24 9
<< metal1 >>
rect -10 -8 -7 19
rect -10 -16 -7 -12
rect -4 16 -1 19
rect -4 12 2 16
rect 27 16 30 19
rect 9 14 13 15
rect -4 0 -1 12
rect 24 12 30 16
rect 6 4 16 7
rect 27 0 30 12
rect -4 -4 2 0
rect 24 -4 30 0
rect -4 -16 -1 -4
rect 9 -16 13 -12
rect 27 -16 30 -4
rect 33 -8 36 19
rect 33 -16 36 -12
<< ntransistor >>
rect 2 9 6 11
<< ptransistor >>
rect 16 9 24 11
<< polycontact >>
rect 9 10 13 14
rect 9 0 13 4
rect -11 -12 -7 -8
rect 33 -12 37 -8
<< ndcontact >>
rect 2 12 6 16
rect 2 4 6 8
<< pdcontact >>
rect 16 12 24 16
rect 16 4 24 8
<< m2contact >>
rect 9 15 13 19
use latch  latch_0
timestamp 1430426212
transform 0 1 2 -1 0 -6
box -6 -2 10 24
<< labels >>
rlabel m2contact 9 15 13 19 5 in
rlabel metal1 -4 16 -1 19 5 GND
rlabel metal1 27 16 30 19 5 Vdd
rlabel metal1 33 16 36 19 6 r_
rlabel metal1 -10 16 -7 19 4 r
rlabel metal1 9 -16 13 -12 1 out
<< end >>
