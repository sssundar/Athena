magic
tech scmos
timestamp 1434148540
<< polysilicon >>
rect 11 1019 21 1021
rect 50 1000 52 1032
rect 107 1017 109 1032
rect 95 1015 109 1017
rect 171 1008 173 1033
rect 81 1006 173 1008
rect 50 998 84 1000
<< metal1 >>
rect 0 989 3 992
rect 7 989 10 1019
rect 14 989 17 1039
rect 45 1032 48 1036
rect 72 1023 75 1038
rect 103 1032 106 1036
rect 130 1023 133 1037
rect 161 1033 169 1037
rect 21 1022 75 1023
rect 25 1020 75 1022
rect 78 1020 133 1023
rect 78 1014 81 1020
rect 21 1011 81 1014
rect 21 989 24 1011
rect 28 989 31 996
rect 70 989 73 992
rect 77 989 80 1004
rect 84 989 87 996
rect 91 989 94 1013
rect 98 989 101 992
rect 105 989 108 992
rect 165 989 168 992
rect 171 989 174 992
rect 200 989 203 992
rect 206 989 209 992
rect 0 867 3 875
rect 7 867 10 875
rect 14 867 17 875
rect 21 867 24 875
rect 28 867 31 875
rect 70 867 73 875
rect 77 867 80 875
rect 84 867 87 875
rect 91 867 94 875
rect 98 867 101 875
rect 105 867 108 875
rect 111 867 114 875
rect 142 867 145 875
rect 165 867 168 880
rect 171 867 174 880
rect 184 867 190 880
rect 200 867 203 880
rect 206 867 209 880
rect 229 867 232 875
rect 0 742 3 750
rect 7 742 10 750
rect 14 742 17 750
rect 21 742 24 750
rect 28 742 31 750
rect 70 742 73 750
rect 77 742 80 750
rect 84 742 87 750
rect 91 742 94 750
rect 98 742 101 750
rect 105 742 108 750
rect 111 742 114 750
rect 142 742 145 750
rect 165 742 168 755
rect 171 742 174 755
rect 184 742 190 755
rect 200 742 203 755
rect 206 742 209 755
rect 229 742 232 750
rect 0 617 3 625
rect 7 617 10 625
rect 14 617 17 625
rect 21 617 24 625
rect 28 617 31 625
rect 70 617 73 625
rect 77 617 80 625
rect 84 617 87 625
rect 91 617 94 625
rect 98 617 101 625
rect 105 617 108 625
rect 111 617 114 625
rect 142 617 145 625
rect 165 617 168 630
rect 171 617 174 630
rect 184 617 190 630
rect 200 617 203 630
rect 206 617 209 630
rect 229 617 232 625
rect 0 492 3 500
rect 7 492 10 500
rect 14 492 17 500
rect 21 492 24 500
rect 28 492 31 500
rect 70 492 73 500
rect 77 492 80 500
rect 84 492 87 500
rect 91 492 94 500
rect 98 492 101 500
rect 105 492 108 500
rect 111 492 114 500
rect 142 492 145 500
rect 165 492 168 505
rect 171 492 174 505
rect 184 492 190 505
rect 200 492 203 505
rect 206 492 209 505
rect 229 492 232 500
rect 0 367 3 375
rect 7 367 10 375
rect 14 367 17 375
rect 21 367 24 375
rect 28 367 31 375
rect 70 367 73 375
rect 77 367 80 375
rect 84 367 87 375
rect 91 367 94 375
rect 98 367 101 375
rect 105 367 108 375
rect 111 367 114 375
rect 142 367 145 375
rect 165 367 168 380
rect 171 367 174 380
rect 184 367 190 380
rect 200 367 203 380
rect 206 367 209 380
rect 229 367 232 375
rect 0 242 3 250
rect 7 242 10 250
rect 14 242 17 250
rect 21 242 24 250
rect 28 242 31 250
rect 70 242 73 250
rect 77 242 80 250
rect 84 242 87 250
rect 91 242 94 250
rect 98 242 101 250
rect 105 242 108 250
rect 111 242 114 250
rect 142 242 145 250
rect 165 242 168 255
rect 171 242 174 255
rect 184 242 190 255
rect 200 242 203 255
rect 206 242 209 255
rect 229 242 232 250
rect 0 117 3 125
rect 7 117 10 125
rect 14 117 17 125
rect 21 117 24 125
rect 28 117 31 125
rect 70 117 73 125
rect 77 117 80 125
rect 84 117 87 125
rect 91 117 94 125
rect 98 117 101 125
rect 105 117 108 125
rect 111 117 114 125
rect 142 117 145 125
rect 165 117 168 130
rect 171 117 174 130
rect 184 117 190 130
rect 200 117 203 130
rect 206 117 209 130
rect 229 117 232 125
rect 105 0 108 3
<< metal2 >>
rect 29 1000 32 1026
<< polycontact >>
rect 48 1032 52 1036
rect 106 1032 110 1036
rect 169 1033 173 1037
rect 7 1019 11 1023
rect 21 1018 25 1022
rect 91 1013 95 1017
rect 77 1004 81 1008
rect 84 996 88 1000
<< m2contact >>
rect 28 996 32 1000
rect 41 988 45 992
rect 41 863 45 867
rect 41 738 45 742
rect 41 613 45 617
rect 41 488 45 492
rect 41 363 45 367
rect 41 238 45 242
rect 41 113 45 117
use fAccumulatorController  fAccumulatorController_0
timestamp 1434090485
transform 1 0 92 0 1 1218
box -91 -192 83 -98
use fcell  f7
timestamp 1434088717
transform 1 0 111 0 1 892
box -111 -17 121 100
use fcell  f6
timestamp 1434088717
transform 1 0 111 0 1 767
box -111 -17 121 100
use fcell  f5
timestamp 1434088717
transform 1 0 111 0 1 642
box -111 -17 121 100
use fcell  f4
timestamp 1434088717
transform 1 0 111 0 1 517
box -111 -17 121 100
use fcell  f3
timestamp 1434088717
transform 1 0 111 0 1 392
box -111 -17 121 100
use fcell  f2
timestamp 1434088717
transform 1 0 111 0 1 267
box -111 -17 121 100
use fcell  f1
timestamp 1434088717
transform 1 0 111 0 1 142
box -111 -17 121 100
use fcell  f0
timestamp 1434088717
transform 1 0 111 0 1 17
box -111 -17 121 100
<< labels >>
rlabel metal1 0 989 3 992 4 phi1
rlabel metal1 7 989 10 992 5 ld
rlabel metal1 14 989 17 992 5 w
rlabel metal1 21 989 24 992 5 r
rlabel metal1 28 989 31 992 5 GND
rlabel metal1 70 989 73 992 5 Vdd
rlabel metal1 77 989 80 992 5 r_
rlabel metal1 84 989 87 992 5 w_
rlabel metal1 91 989 94 992 5 ld_
rlabel metal1 98 989 101 992 5 phi1_
rlabel metal1 105 989 108 992 5 zout
rlabel metal1 165 989 168 992 5 g1_
rlabel metal1 171 989 174 992 5 g2_
rlabel metal1 200 989 203 992 5 g3_
rlabel metal1 206 989 209 992 5 g0_
rlabel metal1 105 0 108 3 1 zin
rlabel m2contact 41 113 45 117 1 bus0
rlabel m2contact 41 238 45 242 1 bus1
rlabel m2contact 41 363 45 367 1 bus2
rlabel m2contact 41 488 45 492 1 bus3
rlabel m2contact 41 613 45 617 1 bus4
rlabel m2contact 41 738 45 742 1 bus5
rlabel m2contact 41 863 45 867 1 bus6
rlabel m2contact 41 988 45 992 5 bus7
<< end >>
