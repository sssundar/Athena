magic
tech scmos
timestamp 1434158785
<< polysilicon >>
rect 115 1036 118 1038
rect 115 1020 117 1036
rect 98 1014 100 1016
<< metal1 >>
rect 118 1040 122 1042
rect 84 1026 87 1034
rect 125 1025 128 1034
rect 111 1021 115 1025
rect 0 985 3 991
rect 7 985 10 991
rect 15 985 18 991
rect 51 985 54 991
rect 57 985 60 991
rect 64 985 67 991
rect 70 988 73 989
rect 77 988 80 989
rect 84 988 87 989
rect 125 988 128 989
rect 131 985 134 988
rect 138 985 141 988
rect 145 985 148 988
rect 188 985 191 988
rect 195 985 198 988
rect 202 985 205 988
rect 0 863 3 875
rect 7 863 10 875
rect 15 863 18 875
rect 51 863 54 875
rect 57 863 60 875
rect 64 863 67 875
rect 70 863 73 875
rect 77 863 80 875
rect 84 863 87 875
rect 125 863 128 875
rect 131 863 134 875
rect 138 863 141 875
rect 145 863 148 875
rect 152 863 155 875
rect 188 863 191 875
rect 195 863 198 875
rect 202 863 205 875
rect 215 863 218 875
rect 222 863 225 875
rect 261 863 264 875
rect 268 863 271 875
rect 0 738 3 750
rect 7 738 10 750
rect 15 738 18 750
rect 51 738 54 750
rect 57 738 60 750
rect 64 738 67 750
rect 70 738 73 750
rect 77 738 80 750
rect 84 738 87 750
rect 125 738 128 750
rect 131 738 134 750
rect 138 738 141 750
rect 145 738 148 750
rect 152 738 155 750
rect 188 738 191 750
rect 195 738 198 750
rect 202 738 205 750
rect 215 738 218 750
rect 222 738 225 750
rect 261 738 264 750
rect 268 738 271 750
rect 0 613 3 625
rect 7 613 10 625
rect 15 613 18 625
rect 51 613 54 625
rect 57 613 60 625
rect 64 613 67 625
rect 70 613 73 625
rect 77 613 80 625
rect 84 613 87 625
rect 125 613 128 625
rect 131 613 134 625
rect 138 613 141 625
rect 145 613 148 625
rect 152 613 155 625
rect 188 613 191 625
rect 195 613 198 625
rect 202 613 205 625
rect 215 613 218 625
rect 222 613 225 625
rect 261 613 264 625
rect 268 613 271 625
rect 0 488 3 500
rect 7 488 10 500
rect 15 488 18 500
rect 51 488 54 500
rect 57 488 60 500
rect 64 488 67 500
rect 70 488 73 500
rect 77 488 80 500
rect 84 488 87 500
rect 125 488 128 500
rect 131 488 134 500
rect 138 488 141 500
rect 145 488 148 500
rect 152 488 155 500
rect 188 488 191 500
rect 195 488 198 500
rect 202 488 205 500
rect 215 488 218 500
rect 222 488 225 500
rect 261 488 264 500
rect 268 488 271 500
rect 0 363 3 375
rect 7 363 10 375
rect 15 363 18 375
rect 51 363 54 375
rect 57 363 60 375
rect 64 363 67 375
rect 70 363 73 375
rect 77 363 80 375
rect 84 363 87 375
rect 125 363 128 375
rect 131 363 134 375
rect 138 363 141 375
rect 145 363 148 375
rect 152 363 155 375
rect 188 363 191 375
rect 195 363 198 375
rect 202 363 205 375
rect 215 363 218 375
rect 222 363 225 375
rect 261 363 264 375
rect 268 363 271 375
rect 0 238 3 250
rect 7 238 10 250
rect 15 238 18 250
rect 51 238 54 250
rect 57 238 60 250
rect 64 238 67 250
rect 70 238 73 250
rect 77 238 80 250
rect 84 238 87 250
rect 125 238 128 250
rect 131 238 134 250
rect 138 238 141 250
rect 145 238 148 250
rect 152 238 155 250
rect 188 238 191 250
rect 195 238 198 250
rect 202 238 205 250
rect 215 238 218 250
rect 222 238 225 250
rect 261 238 264 250
rect 268 238 271 250
rect 0 113 3 125
rect 7 113 10 125
rect 15 113 18 125
rect 51 113 54 125
rect 57 113 60 125
rect 64 113 67 125
rect 70 113 73 125
rect 77 113 80 125
rect 84 113 87 125
rect 125 113 128 125
rect 131 113 134 125
rect 138 113 141 125
rect 145 113 148 125
rect 152 113 155 125
rect 188 113 191 125
rect 195 113 198 125
rect 202 113 205 125
rect 215 113 218 125
rect 222 113 225 125
rect 261 113 264 125
rect 268 113 271 125
<< metal2 >>
rect 29 931 33 935
rect 29 806 33 810
rect 29 681 33 685
rect 29 556 33 560
rect 29 431 33 435
rect 29 306 33 310
rect 29 181 33 185
rect 29 56 33 60
<< polycontact >>
rect 118 1036 122 1040
use pwm_controller  pwm_controller_0
timestamp 1434158785
transform 1 0 0 0 1 0
box 0 991 143 1091
use pwmoutput  pwmoutput_0
timestamp 1433956774
transform -1 0 128 0 1 891
box 0 98 58 135
use pwmcell  pwm7
timestamp 1434158463
transform 1 0 -6 0 1 866
box 6 9 282 122
use pwmcell  pwm6
timestamp 1434158463
transform 1 0 -6 0 1 741
box 6 9 282 122
use pwmcell  pwm5
timestamp 1434158463
transform 1 0 -6 0 1 616
box 6 9 282 122
use pwmcell  pwm4
timestamp 1434158463
transform 1 0 -6 0 1 491
box 6 9 282 122
use pwmcell  pwm3
timestamp 1434158463
transform 1 0 -6 0 1 366
box 6 9 282 122
use pwmcell  pwm2
timestamp 1434158463
transform 1 0 -6 0 1 241
box 6 9 282 122
use pwmcell  pwm1
timestamp 1434158463
transform 1 0 -6 0 1 116
box 6 9 282 122
use pwmcell  pwm0
timestamp 1434158463
transform 1 0 -6 0 1 -9
box 6 9 282 122
<< labels >>
rlabel metal1 0 985 3 988 4 w
rlabel metal1 7 985 10 988 5 r
rlabel metal1 15 985 18 988 5 GND
rlabel metal1 51 985 54 988 5 Vdd
rlabel metal1 57 985 60 988 5 r_
rlabel metal1 64 985 67 988 5 w_
rlabel metal1 111 1021 115 1025 5 pwmout
rlabel polysilicon 98 1014 100 1016 1 pwmoe_
rlabel metal1 131 985 134 988 1 phi1
rlabel metal1 138 985 141 988 1 phi0
rlabel metal1 145 985 148 988 1 reset
rlabel metal1 195 985 198 988 1 phi0_
rlabel metal1 202 985 205 988 1 phi1_
rlabel metal2 29 56 33 60 1 bus0
rlabel metal2 29 181 33 185 1 bus1
rlabel metal2 29 306 33 310 1 bus2
rlabel metal2 29 431 33 435 1 bus3
rlabel metal2 29 556 33 560 1 bus4
rlabel metal2 29 681 33 685 1 bus5
rlabel metal2 29 806 33 810 1 bus6
rlabel metal2 29 931 33 935 1 bus7
<< end >>
