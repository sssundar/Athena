magic
tech scmos
timestamp 1434174869
<< polysilicon >>
rect -60 -86 -48 -84
rect -68 -98 -66 -96
rect -68 -105 -66 -102
rect -68 -109 -67 -105
rect -68 -112 -66 -109
rect -60 -112 -58 -86
rect -46 -89 -41 -87
rect -37 -89 -35 -87
rect -33 -91 -31 -40
rect -22 -87 -20 -40
rect -12 -42 -10 -40
rect -4 -42 -2 -40
rect 0 -42 2 -40
rect 8 -42 10 -40
rect 12 -42 14 -40
rect -12 -48 -10 -46
rect -4 -61 -2 -46
rect -15 -63 -13 -61
rect -5 -63 -2 -61
rect 0 -61 2 -46
rect 8 -51 10 -46
rect 12 -47 14 -46
rect 12 -49 18 -47
rect 8 -53 14 -51
rect 12 -61 14 -53
rect 0 -63 3 -61
rect 11 -63 14 -61
rect 16 -69 18 -49
rect -15 -71 -13 -69
rect -5 -71 -3 -69
rect 1 -71 3 -69
rect 11 -71 18 -69
rect 20 -73 22 -27
rect 28 -42 30 -40
rect 44 -42 46 -40
rect 52 -42 54 -40
rect 56 -42 58 -40
rect 28 -49 30 -46
rect 44 -47 46 -46
rect 29 -53 30 -49
rect 28 -56 30 -53
rect 36 -49 46 -47
rect 52 -48 54 -46
rect 36 -61 38 -49
rect 51 -50 54 -48
rect 36 -63 39 -61
rect 47 -63 49 -61
rect 15 -75 22 -73
rect -29 -89 -27 -87
rect -23 -89 -17 -87
rect -51 -93 -41 -91
rect -37 -93 -35 -91
rect -33 -93 -27 -91
rect -23 -93 -21 -91
rect -53 -109 -51 -94
rect -46 -96 -41 -95
rect -44 -97 -41 -96
rect -37 -97 -35 -95
rect -53 -111 -50 -109
rect -52 -112 -50 -111
rect -44 -112 -42 -97
rect -68 -122 -66 -120
rect -60 -122 -58 -120
rect -52 -122 -50 -120
rect -44 -122 -42 -120
rect -33 -123 -31 -93
rect -19 -119 -17 -89
rect 15 -91 17 -75
rect 28 -86 30 -64
rect 51 -69 53 -50
rect 56 -52 58 -46
rect 37 -71 39 -69
rect 47 -71 53 -69
rect 55 -54 58 -52
rect 55 -69 57 -54
rect 67 -65 69 -40
rect 75 -42 77 -40
rect 75 -49 77 -46
rect 76 -53 77 -49
rect 75 -56 77 -53
rect 67 -67 72 -65
rect 75 -66 77 -64
rect 55 -71 58 -69
rect 66 -71 68 -69
rect 28 -87 31 -86
rect 19 -89 21 -87
rect 25 -89 31 -87
rect -4 -93 21 -91
rect 25 -93 27 -91
rect -4 -96 -2 -93
rect -9 -98 -2 -96
rect -9 -112 -7 -98
rect 12 -101 21 -99
rect 25 -101 27 -99
rect 12 -107 14 -101
rect 0 -109 3 -107
rect 11 -109 14 -107
rect 29 -109 31 -89
rect 70 -91 72 -67
rect 82 -73 83 -71
rect 81 -87 83 -73
rect 74 -89 76 -87
rect 80 -89 86 -87
rect 44 -93 76 -91
rect 80 -93 82 -91
rect 44 -107 46 -93
rect 84 -107 86 -89
rect 33 -109 35 -107
rect 43 -109 46 -107
rect 48 -109 50 -107
rect 58 -109 86 -107
rect -9 -114 -4 -112
rect 28 -111 31 -109
rect -6 -118 -4 -114
rect 31 -117 35 -115
rect 43 -117 45 -115
rect 48 -117 50 -115
rect 58 -117 63 -115
rect 31 -118 33 -117
rect -6 -120 33 -118
rect -33 -125 35 -123
rect 43 -125 45 -123
rect 48 -125 50 -123
rect 58 -125 63 -123
<< ndiffusion >>
rect -69 -102 -68 -98
rect -66 -102 -65 -98
rect -41 -87 -37 -86
rect -41 -91 -37 -89
rect -27 -87 -23 -86
rect -13 -46 -12 -42
rect -10 -46 -9 -42
rect -5 -46 -4 -42
rect -2 -46 0 -42
rect 2 -46 3 -42
rect 7 -46 8 -42
rect 10 -46 12 -42
rect 14 -46 15 -42
rect 27 -46 28 -42
rect 30 -46 31 -42
rect 43 -46 44 -42
rect 46 -46 47 -42
rect 51 -46 52 -42
rect 54 -46 56 -42
rect 58 -46 59 -42
rect -27 -91 -23 -89
rect -41 -95 -37 -93
rect -41 -98 -37 -97
rect -27 -94 -23 -93
rect 21 -87 25 -86
rect 74 -46 75 -42
rect 77 -46 78 -42
rect 21 -91 25 -89
rect 21 -94 25 -93
rect 21 -99 25 -98
rect 21 -102 25 -101
rect 76 -87 80 -86
rect 76 -91 80 -89
rect 76 -94 80 -93
<< pdiffusion >>
rect -13 -61 -5 -60
rect 3 -61 11 -60
rect -13 -64 -5 -63
rect -13 -69 -5 -68
rect 3 -64 11 -63
rect 3 -69 11 -68
rect -13 -72 -5 -71
rect 3 -72 11 -71
rect 27 -64 28 -56
rect 30 -64 31 -56
rect 39 -61 47 -60
rect 39 -64 47 -63
rect -69 -120 -68 -112
rect -66 -120 -65 -112
rect -61 -120 -60 -112
rect -58 -120 -57 -112
rect -53 -120 -52 -112
rect -50 -120 -49 -112
rect -45 -120 -44 -112
rect -42 -120 -41 -112
rect 39 -69 47 -68
rect 74 -64 75 -56
rect 77 -64 78 -56
rect 58 -69 66 -68
rect 39 -72 47 -71
rect 58 -72 66 -71
rect 3 -107 11 -106
rect 35 -107 43 -106
rect 50 -107 58 -106
rect 3 -110 11 -109
rect 35 -110 43 -109
rect 35 -115 43 -114
rect 50 -110 58 -109
rect 50 -115 58 -114
rect 35 -118 43 -117
rect 35 -123 43 -122
rect 50 -118 58 -117
rect 50 -123 58 -122
rect 35 -126 43 -125
rect 50 -126 58 -125
<< metal1 >>
rect -64 -20 42 -17
rect -64 -98 -61 -20
rect -54 -27 19 -24
rect -54 -90 -51 -27
rect -47 -33 35 -30
rect -47 -83 -44 -33
rect -27 -39 26 -36
rect -27 -82 -23 -39
rect -17 -42 -13 -39
rect 3 -42 7 -39
rect 23 -42 26 -39
rect 31 -42 35 -33
rect 39 -36 42 -20
rect 39 -39 89 -36
rect 39 -42 43 -39
rect 59 -42 63 -39
rect 63 -46 70 -42
rect -9 -56 -5 -46
rect 15 -49 19 -46
rect 15 -53 25 -49
rect 15 -56 19 -53
rect 32 -56 35 -46
rect 47 -49 51 -46
rect 47 -53 72 -49
rect -5 -60 3 -56
rect 11 -59 19 -56
rect 47 -60 51 -53
rect 79 -56 82 -46
rect -5 -68 3 -64
rect 23 -72 27 -64
rect 47 -68 58 -64
rect 70 -72 74 -64
rect -5 -76 3 -72
rect 11 -76 39 -72
rect 47 -74 58 -72
rect 47 -76 51 -74
rect 55 -76 58 -74
rect 66 -76 74 -72
rect 78 -69 82 -64
rect 86 -82 89 -39
rect -37 -86 -27 -82
rect -23 -86 21 -82
rect 25 -86 76 -82
rect 80 -86 93 -82
rect -48 -94 -30 -91
rect -48 -96 -44 -94
rect -73 -112 -70 -102
rect -41 -106 -37 -102
rect -63 -109 -37 -106
rect -33 -106 -30 -94
rect -23 -98 21 -94
rect 25 -98 76 -94
rect -33 -109 -4 -106
rect 11 -106 21 -102
rect 25 -106 35 -102
rect 43 -106 50 -102
rect 58 -106 81 -102
rect 89 -105 93 -86
rect -57 -112 -53 -109
rect -41 -112 -37 -109
rect 23 -113 24 -109
rect 43 -114 50 -110
rect 77 -112 81 -106
rect -13 -119 -12 -115
rect -65 -123 -61 -120
rect -49 -123 -45 -120
rect 7 -123 11 -114
rect 67 -118 68 -114
rect 77 -116 90 -112
rect 97 -116 101 -112
rect 43 -122 50 -118
rect -65 -126 11 -123
rect 67 -126 68 -122
rect 7 -129 35 -126
rect 43 -130 50 -126
rect 58 -130 78 -129
rect 54 -131 78 -130
rect 89 -129 92 -127
rect 82 -131 92 -129
rect 54 -132 92 -131
<< metal2 >>
rect 51 -100 55 -78
rect 51 -104 82 -100
rect 23 -113 72 -109
rect 68 -114 72 -113
rect -12 -122 -8 -119
rect -12 -126 68 -122
rect 78 -127 82 -104
<< ntransistor >>
rect -68 -102 -66 -98
rect -41 -89 -37 -87
rect -12 -46 -10 -42
rect -4 -46 -2 -42
rect 0 -46 2 -42
rect 8 -46 10 -42
rect 12 -46 14 -42
rect 28 -46 30 -42
rect 44 -46 46 -42
rect 52 -46 54 -42
rect 56 -46 58 -42
rect -27 -89 -23 -87
rect -41 -93 -37 -91
rect -27 -93 -23 -91
rect -41 -97 -37 -95
rect 75 -46 77 -42
rect 21 -89 25 -87
rect 21 -93 25 -91
rect 21 -101 25 -99
rect 76 -89 80 -87
rect 76 -93 80 -91
<< ptransistor >>
rect -13 -63 -5 -61
rect 3 -63 11 -61
rect -13 -71 -5 -69
rect 3 -71 11 -69
rect 28 -64 30 -56
rect 39 -63 47 -61
rect -68 -120 -66 -112
rect -60 -120 -58 -112
rect -52 -120 -50 -112
rect -44 -120 -42 -112
rect 39 -71 47 -69
rect 75 -64 77 -56
rect 58 -71 66 -69
rect 3 -109 11 -107
rect 35 -109 43 -107
rect 50 -109 58 -107
rect 35 -117 43 -115
rect 50 -117 58 -115
rect 35 -125 43 -123
rect 50 -125 58 -123
<< polycontact >>
rect 19 -27 23 -23
rect -67 -109 -63 -105
rect -48 -87 -44 -83
rect -55 -94 -51 -90
rect 25 -53 29 -49
rect -48 -100 -44 -96
rect 72 -53 76 -49
rect -4 -109 0 -105
rect 78 -73 82 -69
rect 24 -113 28 -109
rect -17 -119 -13 -115
rect 63 -118 67 -114
rect 90 -116 94 -112
rect 63 -126 67 -122
<< ndcontact >>
rect -73 -102 -69 -98
rect -65 -102 -61 -98
rect -41 -86 -37 -82
rect -27 -86 -23 -82
rect -17 -46 -13 -42
rect -9 -46 -5 -42
rect 3 -46 7 -42
rect 15 -46 19 -42
rect 23 -46 27 -42
rect 31 -46 35 -42
rect 39 -46 43 -42
rect 47 -46 51 -42
rect 59 -46 63 -42
rect -41 -102 -37 -98
rect -27 -98 -23 -94
rect 21 -86 25 -82
rect 70 -46 74 -42
rect 78 -46 82 -42
rect 21 -98 25 -94
rect 21 -106 25 -102
rect 76 -86 80 -82
rect 76 -98 80 -94
<< pdcontact >>
rect -13 -60 -5 -56
rect 3 -60 11 -56
rect -13 -68 -5 -64
rect 3 -68 11 -64
rect -13 -76 -5 -72
rect 3 -76 11 -72
rect 23 -64 27 -56
rect 31 -64 35 -56
rect 39 -60 47 -56
rect -73 -120 -69 -112
rect -65 -120 -61 -112
rect -57 -120 -53 -112
rect -49 -120 -45 -112
rect -41 -120 -37 -112
rect 39 -68 47 -64
rect 58 -68 66 -64
rect 70 -64 74 -56
rect 78 -64 82 -56
rect 39 -76 47 -72
rect 58 -76 66 -72
rect 3 -106 11 -102
rect 35 -106 43 -102
rect 50 -106 58 -102
rect 3 -114 11 -110
rect 35 -114 43 -110
rect 50 -114 58 -110
rect 35 -122 43 -118
rect 50 -122 58 -118
rect 35 -130 43 -126
rect 50 -130 58 -126
<< m2contact >>
rect 51 -78 55 -74
rect 19 -113 23 -109
rect -12 -119 -8 -115
rect 68 -118 72 -114
rect 68 -126 72 -122
rect 78 -131 82 -127
use inverter  inverter_0
timestamp 1430424850
transform 1 0 94 0 -1 -98
box -5 5 7 31
<< labels >>
rlabel polysilicon -11 -41 -11 -41 5 ctl4
rlabel polysilicon -3 -41 -3 -41 5 ctl2
rlabel polysilicon 1 -41 1 -41 5 carry
rlabel polysilicon 9 -41 9 -41 5 ctl3
rlabel polysilicon 13 -41 13 -41 3 zero
rlabel metal1 15 -58 15 -58 1 branch_
rlabel metal1 33 -51 33 -51 7 branch
rlabel metal1 49 -51 49 -51 1 shouldinc_
rlabel metal1 80 -51 80 -51 7 shouldinc
rlabel polysilicon 45 -41 45 -41 5 branchinst
rlabel polysilicon 53 -41 53 -41 5 inputinst
rlabel polysilicon 57 -41 57 -41 5 ctl3_
rlabel polysilicon 21 -41 21 -41 5 cnt2
rlabel polysilicon 68 -41 68 -41 5 cnt1
rlabel polysilicon -32 -42 -32 -42 4 cnt0
rlabel polysilicon -21 -42 -21 -42 5 reset_
rlabel polycontact -2 -107 -2 -107 1 phi0
rlabel metal1 -55 -108 -55 -108 1 branch_w_
rlabel ndcontact 21 -106 25 -102 1 inc_w_
rlabel metal1 99 -114 99 -114 7 inc_w
rlabel metal1 -71 -107 -71 -107 3 branch_w
rlabel ndcontact -63 -100 -63 -100 1 GND
rlabel metal1 91 -131 91 -131 1 Vdd
<< end >>
