magic
tech scmos
timestamp 1430475211
<< polysilicon >>
rect -35 83 -33 85
rect -27 83 -25 90
rect -35 48 -33 51
rect -34 44 -33 48
rect -35 41 -33 44
rect -27 41 -25 51
rect -18 45 -9 47
rect -35 23 -33 25
rect -27 23 -25 25
rect -42 8 -40 10
rect -36 8 -26 10
rect -18 8 -16 10
rect -49 -1 -29 1
<< ndiffusion >>
rect -36 25 -35 41
rect -33 25 -27 41
rect -25 25 -24 41
rect -40 10 -36 11
rect -40 7 -36 8
<< pdiffusion >>
rect -36 51 -35 83
rect -33 55 -27 83
rect -33 51 -32 55
rect -28 51 -27 55
rect -25 51 -24 83
rect -26 10 -18 11
rect -26 7 -18 8
<< metal1 >>
rect -30 90 -29 94
rect -40 84 -12 87
rect -40 83 -36 84
rect -24 83 -12 84
rect -16 79 -12 83
rect -39 44 -38 48
rect -31 46 -28 51
rect -24 46 -22 47
rect -31 44 -22 46
rect -31 43 -21 44
rect -24 41 -21 43
rect -38 21 -37 25
rect -24 21 -21 25
rect -46 17 -37 21
rect -52 -2 -49 -1
rect -46 -2 -43 17
rect -40 15 -37 17
rect -32 18 -21 21
rect -32 14 -29 18
rect -15 17 -12 79
rect -14 13 -12 17
rect -18 12 -12 13
rect -36 5 -26 7
rect -36 3 -33 5
rect -29 3 -26 5
rect -15 -2 -12 12
rect -9 -2 -6 44
<< ntransistor >>
rect -35 25 -33 41
rect -27 25 -25 41
rect -40 8 -36 10
<< ptransistor >>
rect -35 51 -33 83
rect -27 51 -25 83
rect -26 8 -18 10
<< polycontact >>
rect -29 90 -25 94
rect -38 44 -34 48
rect -22 44 -18 48
rect -9 44 -5 48
rect -33 10 -29 14
rect -53 -1 -49 3
rect -33 1 -29 5
<< ndcontact >>
rect -40 25 -36 41
rect -24 25 -20 41
rect -40 11 -36 15
rect -40 3 -36 7
<< pdcontact >>
rect -40 51 -36 83
rect -32 51 -28 55
rect -24 51 -20 83
rect -26 11 -18 15
rect -26 3 -18 7
<< m2contact >>
rect -34 90 -30 94
rect -43 44 -39 48
<< psubstratepcontact >>
rect -42 21 -38 25
<< nsubstratencontact >>
rect -20 79 -16 83
rect -18 13 -14 17
<< labels >>
rlabel m2contact -34 90 -30 94 1 regr
rlabel m2contact -43 44 -39 48 1 phi1
rlabel metal1 -15 -2 -12 1 1 Vdd
rlabel metal1 -31 5 -31 5 1 out
rlabel metal1 -9 -2 -6 1 1 r_
rlabel metal1 -46 -2 -43 1 1 GND
rlabel metal1 -52 -2 -49 1 3 r
<< end >>
