magic
tech scmos
timestamp 1434094860
<< polysilicon >>
rect -28 23 -26 25
rect -22 24 -12 25
rect -22 23 -19 24
rect -15 23 -12 24
rect -4 23 -2 25
rect -23 15 -12 17
rect -4 15 -2 17
rect -23 5 -21 15
rect -30 3 -28 5
rect -24 3 -21 5
rect -19 7 -12 9
rect -4 7 -2 9
rect -19 1 -17 7
rect -30 -1 -28 1
rect -24 -1 -17 1
rect -15 -1 -12 1
rect -4 -1 -2 1
rect -15 -3 -13 -1
rect -30 -5 -28 -3
rect -24 -5 -13 -3
rect -30 -9 -28 -7
rect -24 -9 -12 -7
rect -4 -9 -2 -7
<< ndiffusion >>
rect -26 25 -22 26
rect -26 22 -22 23
rect -28 5 -24 6
rect -28 1 -24 3
rect -28 -3 -24 -1
rect -28 -7 -24 -5
rect -28 -10 -24 -9
<< pdiffusion >>
rect -12 25 -4 26
rect -12 22 -4 23
rect -12 17 -4 18
rect -12 14 -4 15
rect -12 9 -4 10
rect -12 6 -4 7
rect -12 1 -4 2
rect -12 -2 -4 -1
rect -12 -7 -4 -6
rect -12 -10 -4 -9
<< metal1 >>
rect -34 22 -31 30
rect -22 27 -12 30
rect -34 18 -26 22
rect -1 22 2 30
rect -34 -10 -31 18
rect -18 14 -15 20
rect -4 18 2 22
rect -18 13 -12 14
rect -28 10 -12 13
rect -18 -2 -15 10
rect -1 6 2 18
rect -4 2 2 6
rect -18 -6 -12 -2
rect -1 -10 2 2
rect -34 -14 -28 -10
rect -4 -14 2 -10
<< ntransistor >>
rect -26 23 -22 25
rect -28 3 -24 5
rect -28 -1 -24 1
rect -28 -5 -24 -3
rect -28 -9 -24 -7
<< ptransistor >>
rect -12 23 -4 25
rect -12 15 -4 17
rect -12 7 -4 9
rect -12 -1 -4 1
rect -12 -9 -4 -7
<< polycontact >>
rect -19 20 -15 24
<< ndcontact >>
rect -26 26 -22 30
rect -26 18 -22 22
rect -28 6 -24 10
rect -28 -14 -24 -10
<< pdcontact >>
rect -12 26 -4 30
rect -12 18 -4 22
rect -12 10 -4 14
rect -12 2 -4 6
rect -12 -6 -4 -2
rect -12 -14 -4 -10
<< labels >>
rlabel metal1 -19 27 -15 30 5 out
rlabel polysilicon -29 4 -29 4 3 a
rlabel polysilicon -29 0 -29 0 3 b
rlabel polysilicon -29 -4 -29 -4 3 c
rlabel polysilicon -29 -8 -29 -8 3 d
<< end >>
