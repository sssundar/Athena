magic
tech scmos
timestamp 1434163595
<< polysilicon >>
rect 22 16 24 26
rect 176 -48 179 -44
<< metal1 >>
rect 57 67 184 71
rect 188 70 336 71
rect 188 67 310 70
rect 57 41 61 67
rect 107 63 111 67
rect 231 57 237 67
rect 314 67 336 70
rect -30 38 -7 41
rect 16 38 61 41
rect -30 -16 -27 38
rect 38 35 44 38
rect 197 29 239 32
rect 197 28 220 29
rect 197 20 200 28
rect 224 28 239 29
rect 288 28 334 31
rect 131 17 200 20
rect -24 13 -4 17
rect 52 15 71 16
rect 321 15 324 28
rect 1826 26 1851 38
rect 52 12 87 15
rect 72 11 79 12
rect 83 11 87 12
rect 321 11 326 15
rect 330 11 336 15
rect 258 -3 262 8
rect 17 -5 40 -3
rect 17 -9 21 -5
rect 25 -9 40 -5
rect 56 -7 105 -3
rect 137 -6 336 -3
rect -30 -20 76 -16
rect 84 -24 90 -21
rect 64 -39 68 -31
rect 87 -36 90 -24
rect 94 -27 97 -14
rect 184 -22 188 -21
rect 269 -21 297 -18
rect 220 -27 224 -21
rect 94 -31 99 -27
rect 294 -33 297 -21
rect 310 -22 317 -21
rect 310 -25 319 -22
rect 311 -27 336 -25
rect 316 -28 336 -27
rect 87 -40 99 -36
rect 212 -39 220 -35
rect 294 -36 301 -33
rect 92 -45 96 -40
rect 92 -49 100 -45
rect 172 -53 175 -48
rect 156 -56 175 -53
rect 78 -65 82 -58
rect 139 -65 142 -63
rect 161 -64 188 -60
rect 78 -66 142 -65
rect 25 -69 142 -66
rect 184 -78 188 -64
rect 212 -78 215 -39
rect 292 -78 296 -48
rect 310 -78 314 -67
rect 333 -78 336 -65
rect 184 -82 336 -78
<< metal2 >>
rect 21 -5 24 -4
rect 21 -65 24 -9
rect 68 -10 71 8
rect 65 -13 71 -10
rect 79 -9 83 8
rect 79 -13 94 -9
rect 64 -27 68 -13
rect 184 -17 188 67
rect 314 66 315 67
rect 220 -17 224 25
rect 188 -21 210 -17
rect 206 -44 210 -21
rect 220 -27 224 -21
rect 310 -17 315 66
rect 326 -9 330 11
rect 326 -13 336 -9
rect 314 -21 315 -17
rect 310 -25 315 -21
rect 206 -48 220 -44
<< polycontact >>
rect 20 12 24 16
rect 68 -39 72 -35
rect 301 -37 305 -33
rect 172 -48 176 -44
<< m2contact >>
rect 184 67 188 71
rect 310 66 314 70
rect 220 25 224 29
rect 68 8 72 12
rect 79 8 83 12
rect 326 11 330 15
rect 21 -9 25 -5
rect 94 -14 98 -10
rect 64 -31 68 -27
rect 184 -21 188 -17
rect 220 -21 224 -17
rect 310 -21 314 -17
rect 21 -69 25 -65
use latchOutputMimic  latchOutputMimic_0
timestamp 1434159590
transform 1 0 6 0 1 22
box -16 -31 17 19
use inv_p32n16  inv_p32n16_0
timestamp 1434159157
transform 1 0 54 0 1 19
box -30 -26 8 16
use nand_p32n32  nand_p32n32_0
timestamp 1434160624
transform 1 0 110 0 1 24
box -23 -31 29 41
use nor_p64n16  nor_p64n16_0
timestamp 1434160163
transform 1 0 250 0 1 23
box -48 -17 38 34
use inv_p8n4  inv_p8n4_0
timestamp 1434159005
transform -1 0 80 0 1 -32
box -6 -26 8 16
use trickyxor2  trickyxor2_0
timestamp 1434144344
transform 1 0 119 0 1 -53
box -20 -11 44 43
use inv_p8n4  inv_p8n4_1
timestamp 1434159005
transform -1 0 186 0 1 -38
box -6 -26 8 16
use trickyxnor2  trickyxnor2_0
timestamp 1434146939
transform 1 0 220 0 1 -72
box 0 4 76 54
use inv_p8n4  inv_p8n4_2
timestamp 1434159005
transform -1 0 312 0 1 -41
box -6 -26 8 16
use PCIncrementorOptimizationLargest_BaseCell  PCIncrementorOptimizationLargest_BaseCell_0
array 0 5 249 0 0 153
timestamp 1434163356
transform 1 0 249 0 1 0
box 87 -82 336 71
<< labels >>
rlabel metal1 -22 15 -22 15 3 chainStart
rlabel metal1 22 39 22 39 1 Vdd
rlabel metal1 25 -6 25 -6 1 GND
rlabel metal1 1843 31 1843 31 1 FINALOUTPUT
<< end >>
