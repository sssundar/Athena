magic
tech scmos
timestamp 1433915764
<< polysilicon >>
rect -2 13 0 15
rect 8 13 14 15
rect -7 9 0 11
rect 8 9 10 11
rect -7 2 -5 9
rect -9 0 -5 2
rect -3 5 0 7
rect 8 5 10 7
rect -9 -19 -7 0
rect -3 -1 -1 5
rect -3 -3 1 -1
rect 0 -7 1 -3
rect -1 -15 1 -7
rect 12 -11 14 13
rect 12 -13 17 -11
rect -1 -17 2 -15
rect 6 -17 8 -15
rect -9 -21 -6 -19
rect -2 -21 0 -19
rect 15 -19 17 -13
rect 8 -21 10 -19
rect 14 -21 17 -19
<< ndiffusion >>
rect 2 -15 6 -14
rect -6 -19 -2 -18
rect 2 -18 6 -17
rect -6 -22 -2 -21
rect 10 -19 14 -18
rect 10 -22 14 -21
<< pdiffusion >>
rect 0 15 8 16
rect 0 11 8 13
rect 0 7 8 9
rect 0 4 8 5
<< metal1 >>
rect 3 -10 6 0
rect -6 -14 2 -11
rect 6 -14 14 -11
rect -2 -25 10 -22
<< ntransistor >>
rect 2 -17 6 -15
rect -6 -21 -2 -19
rect 10 -21 14 -19
<< ptransistor >>
rect 0 13 8 15
rect 0 9 8 11
rect 0 5 8 7
<< polycontact >>
rect -4 -7 0 -3
<< ndcontact >>
rect -6 -18 -2 -14
rect 2 -14 6 -10
rect 2 -22 6 -18
rect 10 -18 14 -14
rect -6 -26 -2 -22
rect 10 -26 14 -22
<< pdcontact >>
rect 0 16 8 20
rect 0 0 8 4
<< labels >>
rlabel polycontact -2 -5 -2 -5 1 c
rlabel polysilicon -6 10 -6 10 3 b
rlabel polysilicon -1 14 -1 14 1 a
rlabel pdcontact 4 18 4 18 5 Vdd
rlabel metal1 4 -24 4 -24 1 GND
rlabel metal1 5 -5 5 -5 1 out
<< end >>
