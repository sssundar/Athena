magic
tech scmos
timestamp 1434159590
<< polysilicon >>
rect -16 15 -13 17
rect -16 -20 -14 15
rect -7 8 -5 10
rect 3 8 11 10
rect -8 4 -5 6
rect 3 4 5 6
rect -8 -5 -6 4
rect -8 -16 -6 -9
rect -8 -18 -3 -16
rect 1 -18 3 -16
rect -16 -22 -3 -20
rect 1 -22 3 -20
rect 9 -27 11 8
<< ndiffusion >>
rect -3 -16 1 -15
rect -3 -20 1 -18
rect -3 -23 1 -22
<< pdiffusion >>
rect -5 10 3 11
rect -5 6 3 8
rect -5 3 3 4
<< metal1 >>
rect -9 16 -5 19
rect 3 16 10 19
rect -3 -5 1 -1
rect -3 -9 17 -5
rect -3 -11 1 -9
rect 1 -31 7 -27
<< ntransistor >>
rect -3 -18 1 -16
rect -3 -22 1 -20
<< ptransistor >>
rect -5 8 3 10
rect -5 4 3 6
<< polycontact >>
rect -13 15 -9 19
rect -10 -9 -6 -5
rect 7 -31 11 -27
<< ndcontact >>
rect -3 -15 1 -11
rect -3 -27 1 -23
<< pdcontact >>
rect -5 11 3 15
rect -5 -1 3 3
<< psubstratepcontact >>
rect -3 -31 1 -27
<< nsubstratencontact >>
rect -5 15 3 19
<< labels >>
rlabel polycontact -8 -7 -8 -7 1 flip0to1
rlabel metal1 15 -7 15 -7 7 latchReadMimic
<< end >>
