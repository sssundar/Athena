magic
tech scmos
timestamp 1430424850
<< polysilicon >>
rect 0 29 2 31
rect 0 11 2 21
rect 0 5 2 7
<< ndiffusion >>
rect -1 7 0 11
rect 2 7 3 11
<< pdiffusion >>
rect -1 21 0 29
rect 2 21 3 29
<< metal1 >>
rect 3 11 7 21
<< ntransistor >>
rect 0 7 2 11
<< ptransistor >>
rect 0 21 2 29
<< ndcontact >>
rect -5 7 -1 11
rect 3 7 7 11
<< pdcontact >>
rect -5 21 -1 29
rect 3 21 7 29
<< labels >>
rlabel metal1 5 16 5 16 7 out
<< end >>
