magic
tech scmos
timestamp 1434160018
<< polysilicon >>
rect 0 23 2 25
rect 18 23 28 25
rect 0 19 2 21
rect 18 19 24 21
rect 22 13 24 19
rect 1 11 24 13
rect 1 7 3 11
rect 26 8 28 23
rect -7 5 3 7
rect 1 1 3 5
rect 18 6 28 8
rect 18 4 19 6
rect 17 1 19 4
rect 1 -5 3 -3
rect 17 -5 19 -3
<< ndiffusion >>
rect 0 -3 1 1
rect 3 -3 4 1
rect 16 -3 17 1
rect 19 -3 20 1
<< pdiffusion >>
rect 2 25 18 26
rect 2 21 18 23
rect 2 18 18 19
<< metal1 >>
rect -4 14 2 18
rect 18 14 24 18
rect -4 1 -1 14
rect 21 8 24 14
rect 8 4 14 7
rect 21 5 38 8
rect 8 1 12 4
rect 21 1 24 5
<< ntransistor >>
rect 1 -3 3 1
rect 17 -3 19 1
<< ptransistor >>
rect 2 23 18 25
rect 2 19 18 21
<< polycontact >>
rect -11 5 -7 9
rect 14 4 18 8
<< ndcontact >>
rect -4 -3 0 1
rect 4 -3 8 1
rect 12 -3 16 1
rect 20 -3 24 1
<< pdcontact >>
rect 2 26 18 30
rect 2 14 18 18
<< psubstratepcontact >>
rect 8 -3 12 1
<< nsubstratencontact >>
rect 2 30 18 34
<< labels >>
rlabel polycontact -9 7 -9 7 3 cin
rlabel metal1 36 6 36 6 7 cout
<< end >>
