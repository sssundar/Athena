magic
tech scmos
timestamp 1434159157
<< polysilicon >>
rect -30 5 -28 7
rect 4 5 8 7
rect 6 -15 8 5
rect -16 -17 -14 -15
rect 2 -17 8 -15
<< ndiffusion >>
rect -14 -15 2 -14
rect -14 -18 2 -17
<< pdiffusion >>
rect -28 7 4 8
rect -28 4 4 5
<< metal1 >>
rect -2 -10 2 0
<< ntransistor >>
rect -14 -17 2 -15
<< ptransistor >>
rect -28 5 4 7
<< ndcontact >>
rect -14 -14 2 -10
rect -14 -22 2 -18
<< pdcontact >>
rect -28 8 4 12
rect -28 0 4 4
<< psubstratepcontact >>
rect -14 -26 2 -22
<< nsubstratencontact >>
rect -28 12 4 16
<< end >>
