magic
tech scmos
timestamp 1433960711
<< polysilicon >>
rect 14 21 16 23
rect -7 9 4 11
rect 32 9 41 11
rect -1 -5 1 9
rect 3 -1 5 7
rect 3 -3 6 -1
rect 10 -3 20 -1
rect 28 -3 30 -1
rect -1 -7 6 -5
rect 10 -7 16 -5
rect 14 -9 16 -7
rect 14 -11 20 -9
rect 28 -11 30 -9
rect 30 -27 41 -25
rect -7 -35 13 -33
<< ndiffusion >>
rect 6 -1 10 0
rect 6 -5 10 -3
rect 6 -8 10 -7
<< pdiffusion >>
rect 20 -1 28 0
rect 20 -4 28 -3
rect 20 -9 28 -8
rect 20 -12 28 -11
<< metal1 >>
rect -11 12 -8 31
rect -4 28 -1 31
rect 35 28 38 31
rect -4 24 6 28
rect 28 24 38 28
rect -4 4 -1 24
rect 13 4 17 12
rect 35 4 38 24
rect 42 12 45 31
rect -4 0 6 4
rect 28 0 38 4
rect -4 -20 -1 0
rect 13 -8 20 -4
rect 10 -12 17 -8
rect 35 -12 38 0
rect -4 -24 6 -20
rect 13 -21 17 -12
rect 28 -16 38 -12
rect 35 -20 38 -16
rect -4 -35 -1 -24
rect 28 -24 38 -20
rect 35 -35 38 -24
rect 42 -35 45 -28
<< ntransistor >>
rect 6 -3 10 -1
rect 6 -7 10 -5
<< ptransistor >>
rect 20 -3 28 -1
rect 20 -11 28 -9
<< polycontact >>
rect -11 8 -7 12
rect 41 8 45 12
rect 13 -25 17 -21
rect 41 -28 45 -24
rect -11 -35 -7 -31
rect 13 -35 17 -31
<< ndcontact >>
rect 6 0 10 4
rect 6 -12 10 -8
<< pdcontact >>
rect 20 0 28 4
rect 20 -8 28 -4
rect 20 -16 28 -12
<< m2contact >>
rect 13 0 17 4
use xor  xor_0
timestamp 1433978507
transform 1 0 6 0 1 0
box -6 0 28 31
use inverter  inverter_0
timestamp 1430424850
transform 0 1 -1 -1 0 -25
box -5 5 7 31
<< labels >>
rlabel polycontact -11 -35 -8 -32 2 cout
rlabel m2contact 13 0 17 4 1 s
rlabel metal1 -11 28 -8 31 4 cin
rlabel metal1 42 28 45 31 6 cin_
rlabel metal1 35 28 38 31 5 Vdd
rlabel metal1 -4 28 -1 31 5 GND
rlabel polysilicon 14 21 16 23 1 a_
rlabel polysilicon 3 5 5 7 1 a
rlabel metal1 42 -35 45 -32 8 cout_
<< end >>
