magic
tech scmos
timestamp 1430467387
<< polysilicon >>
rect -45 39 3 40
rect -41 38 3 39
rect -29 31 -4 32
rect -61 28 -31 30
rect -61 5 -59 28
rect -27 30 0 31
rect -7 21 0 23
rect 26 21 46 23
rect -56 15 -51 16
rect -52 14 -51 15
rect -25 15 -20 16
rect -25 14 -24 15
rect 26 10 33 11
rect 26 9 35 10
rect -13 7 -4 9
rect -61 3 -49 5
rect -6 5 0 7
rect 26 5 40 7
rect -26 2 -8 4
rect -10 -1 -8 2
rect -10 -3 10 -1
rect -30 -6 -15 -4
rect -56 -20 -51 -19
rect -52 -21 -51 -20
rect -25 -20 -20 -19
rect -25 -21 -24 -20
rect -17 -36 -15 -6
rect -17 -38 27 -36
<< metal1 >>
rect -56 15 -53 42
rect -45 25 -41 35
rect -38 23 -35 42
rect -31 25 -27 27
rect -23 15 -20 42
rect -56 -20 -53 11
rect -37 6 -33 10
rect -49 -6 -45 2
rect -42 2 -30 6
rect -42 -12 -38 2
rect -34 -10 -30 -6
rect -23 -20 -20 11
rect -56 -39 -53 -24
rect -38 -39 -35 -26
rect -23 -39 -20 -24
rect -17 11 -14 42
rect -10 24 -7 42
rect -17 -39 -14 7
rect -10 -39 -7 20
rect -4 35 -1 42
rect 27 39 30 42
rect 7 36 30 39
rect -4 16 -1 31
rect -4 12 6 16
rect 27 15 30 36
rect -4 -23 -1 12
rect 9 0 12 14
rect 24 12 30 15
rect 9 -4 10 0
rect 27 -4 30 12
rect 33 14 37 15
rect 40 8 43 42
rect 47 24 50 42
rect 9 -8 12 -4
rect 27 -7 35 -4
rect 32 -23 35 -7
rect -4 -27 2 -23
rect 27 -27 35 -23
rect -4 -39 -1 -27
rect 27 -34 30 -27
rect 27 -39 30 -38
rect 40 -39 43 4
rect 47 -39 50 20
<< polycontact >>
rect -45 35 -41 39
rect 3 36 7 40
rect -4 31 0 35
rect -31 27 -27 31
rect -38 19 -34 23
rect -11 20 -7 24
rect 46 20 50 24
rect -56 11 -52 15
rect -24 11 -20 15
rect 9 14 13 18
rect -17 7 -13 11
rect 33 10 37 14
rect -49 2 -45 6
rect -30 2 -26 6
rect 40 4 44 8
rect -34 -6 -30 -2
rect 10 -4 14 0
rect -42 -16 -38 -12
rect -56 -24 -52 -20
rect -24 -24 -20 -20
rect 27 -38 31 -34
<< m2contact >>
rect 9 26 13 30
rect 33 15 37 19
<< psubstratepcontact >>
rect -49 -10 -45 -6
use latch  latch_2
timestamp 1430426212
transform 0 -1 -27 -1 0 19
box -6 -2 10 24
use latch  latch_1
timestamp 1430426212
transform 0 1 2 1 0 18
box -6 -2 10 24
use latch  latch_0
timestamp 1430426212
transform 0 1 2 -1 0 10
box -6 -2 10 24
use latch  latch_3
timestamp 1430426212
transform 0 1 -49 -1 0 -16
box -6 -2 10 24
use staticizer  staticizer_0
timestamp 1430428783
transform 0 1 -2 -1 0 -23
box -19 2 12 32
<< labels >>
rlabel m2contact 33 15 37 19 1 in
rlabel m2contact 9 26 13 30 5 out
rlabel metal1 -38 -39 -35 -36 1 sout
rlabel metal1 -38 39 -35 42 5 sin
rlabel metal1 -56 39 -53 42 5 shift_
rlabel metal1 -23 39 -20 42 5 shift
rlabel metal1 -17 39 -14 42 5 w
rlabel metal1 -10 39 -7 42 5 r
rlabel metal1 -4 39 -1 42 5 GND
rlabel metal1 27 39 30 42 5 VDD
rlabel metal1 40 39 43 42 5 w_
rlabel metal1 47 39 50 42 6 r_
<< end >>
