magic
tech scmos
timestamp 1432009782
<< polysilicon >>
rect 411 19 418 21
rect 422 19 426 21
rect 430 19 434 21
rect 438 19 442 21
rect 446 19 450 21
rect 454 19 458 21
rect 462 19 466 21
rect 470 19 474 21
rect 478 19 482 21
rect 486 19 490 21
rect 494 19 506 21
rect 510 19 514 21
rect 518 19 522 21
rect 526 19 530 21
rect 534 19 538 21
rect 542 19 546 21
rect 550 19 554 21
rect 558 19 565 21
rect 30 12 36 17
rect 30 11 31 12
rect 35 11 36 12
rect 38 12 44 17
rect 38 11 39 12
rect 43 11 44 12
rect 46 12 52 17
rect 46 11 47 12
rect 51 11 52 12
rect 54 12 60 17
rect 54 11 55 12
rect 59 11 60 12
rect 62 12 68 17
rect 62 11 63 12
rect 67 11 68 12
rect 70 12 76 17
rect 70 11 71 12
rect 75 11 76 12
rect 78 12 84 17
rect 78 11 79 12
rect 83 11 84 12
rect 86 12 92 17
rect 86 11 87 12
rect 91 11 92 12
rect 94 12 100 17
rect 94 11 95 12
rect 99 11 100 12
rect 102 12 108 17
rect 102 11 103 12
rect 107 11 108 12
rect 110 12 116 17
rect 110 11 111 12
rect 115 11 116 12
rect 118 12 124 17
rect 118 11 119 12
rect 123 11 124 12
rect 126 12 132 17
rect 126 11 127 12
rect 131 11 132 12
rect 134 12 140 17
rect 134 11 135 12
rect 139 11 140 12
rect 142 12 148 17
rect 142 11 143 12
rect 147 11 148 12
rect 150 12 156 17
rect 150 11 151 12
rect 155 11 156 12
rect 158 12 164 17
rect 158 11 159 12
rect 163 11 164 12
rect 166 12 172 17
rect 166 11 167 12
rect 171 11 172 12
rect 174 12 180 17
rect 174 11 175 12
rect 179 11 180 12
rect 182 12 188 17
rect 182 11 183 12
rect 187 11 188 12
rect 190 12 196 17
rect 190 11 191 12
rect 195 11 196 12
rect 198 12 204 17
rect 198 11 199 12
rect 203 11 204 12
rect 9 -2 11 3
rect 9 -10 11 -6
rect 9 -18 11 -14
rect 9 -26 11 -22
rect 9 -34 11 -30
rect 9 -42 11 -38
rect 9 -50 11 -46
rect 9 -58 11 -54
rect 9 -66 11 -62
rect 9 -74 11 -70
rect 9 -82 11 -78
rect 9 -90 11 -86
rect 9 -98 11 -94
rect 9 -106 11 -102
rect 9 -130 11 -110
rect 9 -138 11 -134
rect 9 -146 11 -142
rect 9 -154 11 -150
rect 9 -162 11 -158
rect 9 -170 11 -166
rect 9 -178 11 -174
rect 9 -186 11 -182
rect 9 -194 11 -190
rect 9 -202 11 -198
rect 9 -210 11 -206
rect 9 -218 11 -214
rect 9 -226 11 -222
rect 9 -234 11 -230
rect 9 -258 11 -238
rect 9 -266 11 -262
rect 9 -274 11 -270
rect 9 -282 11 -278
rect 9 -290 11 -286
rect 9 -298 11 -294
rect 9 -306 11 -302
rect 9 -314 11 -310
rect 9 -322 11 -318
rect 9 -330 11 -326
rect 9 -338 11 -334
rect 9 -346 11 -342
rect 9 -354 11 -350
rect 9 -363 11 -358
rect 31 -368 33 8
rect 39 -2 41 8
rect 39 -10 41 -6
rect 39 -18 41 -14
rect 47 -18 49 8
rect 55 -10 57 8
rect 63 -10 65 8
rect 39 -26 41 -22
rect 39 -34 41 -30
rect 39 -42 41 -38
rect 39 -50 41 -46
rect 39 -58 41 -54
rect 39 -66 41 -62
rect 39 -74 41 -70
rect 39 -82 41 -78
rect 39 -154 41 -86
rect 39 -162 41 -158
rect 47 -162 49 -22
rect 55 -34 57 -14
rect 39 -170 41 -166
rect 39 -202 41 -174
rect 39 -218 41 -206
rect 39 -226 41 -222
rect 39 -258 41 -230
rect 39 -274 41 -262
rect 39 -282 41 -278
rect 39 -290 41 -286
rect 39 -322 41 -294
rect 39 -330 41 -326
rect 39 -338 41 -334
rect 39 -346 41 -342
rect 39 -354 41 -350
rect 39 -368 41 -358
rect 47 -368 49 -166
rect 55 -368 57 -38
rect 63 -154 65 -14
rect 71 -18 73 8
rect 63 -368 65 -158
rect 71 -368 73 -22
rect 79 -26 81 8
rect 79 -368 81 -30
rect 87 -58 89 8
rect 95 -50 97 8
rect 103 -2 105 8
rect 111 -2 113 8
rect 87 -74 89 -62
rect 87 -368 89 -78
rect 95 -368 97 -54
rect 103 -368 105 -6
rect 111 -368 113 -6
rect 119 -42 121 8
rect 127 -2 129 8
rect 127 -42 129 -6
rect 135 -10 137 8
rect 135 -18 137 -14
rect 135 -34 137 -22
rect 143 -34 145 8
rect 151 -2 153 8
rect 151 -10 153 -6
rect 151 -26 153 -14
rect 119 -368 121 -46
rect 127 -50 129 -46
rect 127 -58 129 -54
rect 127 -74 129 -62
rect 135 -66 137 -38
rect 143 -66 145 -38
rect 151 -42 153 -30
rect 151 -50 153 -46
rect 151 -58 153 -54
rect 159 -58 161 8
rect 167 -2 169 8
rect 167 -10 169 -6
rect 167 -18 169 -14
rect 167 -26 169 -22
rect 175 -26 177 8
rect 183 -2 185 8
rect 183 -10 185 -6
rect 167 -34 169 -30
rect 167 -42 169 -38
rect 167 -50 169 -46
rect 127 -82 129 -78
rect 127 -90 129 -86
rect 127 -138 129 -94
rect 135 -98 137 -70
rect 143 -98 145 -70
rect 151 -74 153 -62
rect 159 -66 161 -62
rect 151 -82 153 -78
rect 159 -82 161 -70
rect 167 -74 169 -54
rect 175 -66 177 -30
rect 183 -34 185 -14
rect 191 -26 193 8
rect 199 -2 201 8
rect 220 5 222 7
rect 226 5 236 7
rect 240 5 243 7
rect 247 5 276 7
rect 280 5 290 7
rect 294 5 296 7
rect 212 -3 222 -1
rect 226 -3 247 -1
rect 251 -3 253 -1
rect 303 3 309 4
rect 303 -1 308 3
rect 312 0 343 2
rect 363 0 373 2
rect 383 0 385 2
rect 265 -3 268 -1
rect 272 -3 290 -1
rect 294 -3 296 -1
rect 303 -2 309 -1
rect 199 -10 201 -6
rect 212 -12 214 -3
rect 220 -11 222 -9
rect 226 -11 236 -9
rect 240 -11 243 -9
rect 199 -18 201 -14
rect 303 -5 309 -4
rect 413 -3 418 -1
rect 422 -3 450 -1
rect 454 -3 570 -1
rect 303 -9 308 -5
rect 312 -8 313 -6
rect 333 -8 393 -6
rect 403 -8 405 -6
rect 247 -11 276 -9
rect 280 -11 290 -9
rect 294 -11 296 -9
rect 303 -10 309 -9
rect 212 -19 222 -17
rect 226 -19 247 -17
rect 251 -19 253 -17
rect 303 -13 309 -12
rect 303 -17 308 -13
rect 413 -11 418 -9
rect 422 -11 426 -9
rect 430 -11 434 -9
rect 438 -11 570 -9
rect 312 -16 343 -14
rect 363 -16 373 -14
rect 383 -16 385 -14
rect 265 -19 268 -17
rect 272 -19 290 -17
rect 294 -19 296 -17
rect 303 -18 309 -17
rect 183 -58 185 -38
rect 175 -74 177 -70
rect 151 -90 153 -86
rect 159 -90 161 -86
rect 135 -106 137 -102
rect 143 -106 145 -102
rect 135 -130 137 -110
rect 143 -130 145 -110
rect 127 -146 129 -142
rect 127 -170 129 -150
rect 135 -154 137 -134
rect 135 -162 137 -158
rect 127 -202 129 -174
rect 135 -178 137 -166
rect 135 -186 137 -182
rect 143 -186 145 -134
rect 151 -138 153 -94
rect 159 -98 161 -94
rect 159 -106 161 -102
rect 159 -130 161 -110
rect 151 -146 153 -142
rect 151 -170 153 -150
rect 159 -154 161 -134
rect 167 -138 169 -78
rect 175 -106 177 -78
rect 183 -82 185 -62
rect 191 -66 193 -30
rect 199 -42 201 -22
rect 212 -28 214 -19
rect 220 -27 222 -25
rect 226 -27 236 -25
rect 240 -27 243 -25
rect 303 -21 309 -20
rect 413 -19 418 -17
rect 422 -19 570 -17
rect 303 -25 308 -21
rect 312 -24 313 -22
rect 333 -24 393 -22
rect 403 -24 405 -22
rect 247 -27 276 -25
rect 280 -27 290 -25
rect 294 -27 296 -25
rect 303 -26 309 -25
rect 212 -35 222 -33
rect 226 -35 247 -33
rect 251 -35 253 -33
rect 303 -29 309 -28
rect 303 -33 308 -29
rect 413 -27 434 -25
rect 438 -27 570 -25
rect 312 -32 343 -30
rect 363 -32 373 -30
rect 383 -32 385 -30
rect 265 -35 268 -33
rect 272 -35 290 -33
rect 294 -35 296 -33
rect 303 -34 309 -33
rect 212 -44 214 -35
rect 220 -43 222 -41
rect 226 -43 236 -41
rect 240 -43 243 -41
rect 199 -50 201 -46
rect 303 -37 309 -36
rect 413 -35 418 -33
rect 422 -35 570 -33
rect 303 -41 308 -37
rect 312 -40 313 -38
rect 333 -40 393 -38
rect 403 -40 405 -38
rect 247 -43 276 -41
rect 280 -43 290 -41
rect 294 -43 296 -41
rect 303 -42 309 -41
rect 212 -51 222 -49
rect 226 -51 247 -49
rect 251 -51 253 -49
rect 303 -45 309 -44
rect 303 -49 308 -45
rect 413 -43 426 -41
rect 430 -43 450 -41
rect 454 -43 570 -41
rect 312 -48 343 -46
rect 363 -48 373 -46
rect 383 -48 385 -46
rect 265 -51 268 -49
rect 272 -51 290 -49
rect 294 -51 296 -49
rect 303 -50 309 -49
rect 183 -90 185 -86
rect 191 -90 193 -70
rect 199 -82 201 -54
rect 212 -60 214 -51
rect 220 -59 222 -57
rect 226 -59 236 -57
rect 240 -59 243 -57
rect 303 -53 309 -52
rect 413 -51 426 -49
rect 430 -51 450 -49
rect 454 -51 570 -49
rect 303 -57 308 -53
rect 312 -56 313 -54
rect 333 -56 393 -54
rect 403 -56 405 -54
rect 247 -59 276 -57
rect 280 -59 290 -57
rect 294 -59 296 -57
rect 303 -58 309 -57
rect 212 -67 222 -65
rect 226 -67 247 -65
rect 251 -67 253 -65
rect 303 -61 309 -60
rect 303 -65 308 -61
rect 413 -59 418 -57
rect 422 -59 434 -57
rect 438 -59 450 -57
rect 454 -59 570 -57
rect 312 -64 343 -62
rect 363 -64 373 -62
rect 383 -64 385 -62
rect 265 -67 268 -65
rect 272 -67 290 -65
rect 294 -67 296 -65
rect 303 -66 309 -65
rect 212 -76 214 -67
rect 220 -75 222 -73
rect 226 -75 236 -73
rect 240 -75 243 -73
rect 303 -69 309 -68
rect 413 -67 450 -65
rect 454 -67 570 -65
rect 303 -73 308 -69
rect 312 -72 313 -70
rect 333 -72 393 -70
rect 403 -72 405 -70
rect 247 -75 276 -73
rect 280 -75 290 -73
rect 294 -75 296 -73
rect 303 -74 309 -73
rect 212 -83 222 -81
rect 226 -83 247 -81
rect 251 -83 253 -81
rect 303 -77 309 -76
rect 303 -81 308 -77
rect 413 -75 418 -73
rect 422 -75 426 -73
rect 430 -75 570 -73
rect 312 -80 343 -78
rect 363 -80 373 -78
rect 383 -80 385 -78
rect 265 -83 268 -81
rect 272 -83 290 -81
rect 294 -83 296 -81
rect 303 -82 309 -81
rect 183 -98 185 -94
rect 191 -98 193 -94
rect 175 -130 177 -110
rect 175 -138 177 -134
rect 167 -146 169 -142
rect 151 -178 153 -174
rect 159 -178 161 -158
rect 167 -170 169 -150
rect 135 -194 137 -190
rect 143 -194 145 -190
rect 127 -306 129 -206
rect 135 -210 137 -198
rect 135 -218 137 -214
rect 143 -218 145 -198
rect 151 -202 153 -182
rect 151 -210 153 -206
rect 135 -226 137 -222
rect 135 -234 137 -230
rect 135 -266 137 -238
rect 135 -282 137 -270
rect 135 -290 137 -286
rect 135 -298 137 -294
rect 143 -298 145 -222
rect 151 -226 153 -214
rect 159 -226 161 -182
rect 167 -186 169 -174
rect 175 -178 177 -142
rect 183 -146 185 -102
rect 191 -106 193 -102
rect 191 -138 193 -110
rect 199 -130 201 -86
rect 212 -92 214 -83
rect 220 -91 222 -89
rect 226 -91 236 -89
rect 240 -91 243 -89
rect 303 -85 309 -84
rect 413 -83 434 -81
rect 438 -83 450 -81
rect 454 -83 570 -81
rect 303 -89 308 -85
rect 312 -88 313 -86
rect 333 -88 393 -86
rect 403 -88 405 -86
rect 247 -91 276 -89
rect 280 -91 290 -89
rect 294 -91 296 -89
rect 303 -90 309 -89
rect 212 -99 222 -97
rect 226 -99 247 -97
rect 251 -99 253 -97
rect 303 -93 309 -92
rect 303 -97 308 -93
rect 413 -91 474 -89
rect 478 -91 490 -89
rect 494 -91 570 -89
rect 312 -96 343 -94
rect 363 -96 373 -94
rect 383 -96 385 -94
rect 265 -99 268 -97
rect 272 -99 290 -97
rect 294 -99 296 -97
rect 303 -98 309 -97
rect 212 -108 214 -99
rect 303 -101 309 -100
rect 413 -99 514 -97
rect 518 -99 570 -97
rect 303 -105 308 -101
rect 312 -104 313 -102
rect 333 -104 393 -102
rect 403 -104 405 -102
rect 303 -106 309 -105
rect 413 -107 546 -105
rect 550 -107 570 -105
rect 220 -123 222 -121
rect 226 -123 236 -121
rect 240 -123 243 -121
rect 247 -123 276 -121
rect 280 -123 290 -121
rect 294 -123 296 -121
rect 212 -131 222 -129
rect 226 -131 247 -129
rect 251 -131 253 -129
rect 303 -125 309 -124
rect 303 -129 308 -125
rect 312 -128 343 -126
rect 363 -128 373 -126
rect 383 -128 385 -126
rect 265 -131 268 -129
rect 272 -131 290 -129
rect 294 -131 296 -129
rect 303 -130 309 -129
rect 191 -146 193 -142
rect 183 -162 185 -150
rect 191 -162 193 -150
rect 199 -154 201 -134
rect 212 -140 214 -131
rect 220 -139 222 -137
rect 226 -139 236 -137
rect 240 -139 243 -137
rect 303 -133 309 -132
rect 413 -131 530 -129
rect 534 -131 570 -129
rect 303 -137 308 -133
rect 312 -136 313 -134
rect 333 -136 393 -134
rect 403 -136 405 -134
rect 247 -139 276 -137
rect 280 -139 290 -137
rect 294 -139 296 -137
rect 303 -138 309 -137
rect 212 -147 222 -145
rect 226 -147 247 -145
rect 251 -147 253 -145
rect 303 -141 309 -140
rect 303 -145 308 -141
rect 413 -139 466 -137
rect 470 -139 522 -137
rect 526 -139 570 -137
rect 312 -144 343 -142
rect 363 -144 373 -142
rect 383 -144 385 -142
rect 265 -147 268 -145
rect 272 -147 290 -145
rect 294 -147 296 -145
rect 303 -146 309 -145
rect 212 -156 214 -147
rect 220 -155 222 -153
rect 226 -155 236 -153
rect 240 -155 243 -153
rect 183 -170 185 -166
rect 191 -170 193 -166
rect 175 -186 177 -182
rect 167 -194 169 -190
rect 175 -194 177 -190
rect 167 -202 169 -198
rect 175 -202 177 -198
rect 167 -210 169 -206
rect 175 -210 177 -206
rect 151 -234 153 -230
rect 151 -258 153 -238
rect 151 -266 153 -262
rect 151 -274 153 -270
rect 127 -368 129 -310
rect 135 -314 137 -302
rect 135 -322 137 -318
rect 143 -322 145 -302
rect 151 -306 153 -278
rect 159 -282 161 -230
rect 167 -234 169 -214
rect 175 -218 177 -214
rect 175 -226 177 -222
rect 167 -258 169 -238
rect 167 -266 169 -262
rect 175 -266 177 -230
rect 183 -234 185 -174
rect 191 -194 193 -174
rect 199 -178 201 -158
rect 303 -149 309 -148
rect 413 -147 506 -145
rect 510 -147 530 -145
rect 534 -147 570 -145
rect 303 -153 308 -149
rect 312 -152 313 -150
rect 333 -152 393 -150
rect 403 -152 405 -150
rect 247 -155 276 -153
rect 280 -155 290 -153
rect 294 -155 296 -153
rect 303 -154 309 -153
rect 212 -163 222 -161
rect 226 -163 247 -161
rect 251 -163 253 -161
rect 303 -157 309 -156
rect 303 -161 308 -157
rect 413 -155 418 -153
rect 422 -155 570 -153
rect 312 -160 343 -158
rect 363 -160 373 -158
rect 383 -160 385 -158
rect 265 -163 268 -161
rect 272 -163 290 -161
rect 294 -163 296 -161
rect 303 -162 309 -161
rect 212 -172 214 -163
rect 220 -171 222 -169
rect 226 -171 236 -169
rect 240 -171 243 -169
rect 303 -165 309 -164
rect 413 -163 426 -161
rect 430 -163 570 -161
rect 303 -169 308 -165
rect 312 -168 313 -166
rect 333 -168 393 -166
rect 403 -168 405 -166
rect 247 -171 276 -169
rect 280 -171 290 -169
rect 294 -171 296 -169
rect 303 -170 309 -169
rect 212 -179 222 -177
rect 226 -179 247 -177
rect 251 -179 253 -177
rect 303 -173 309 -172
rect 303 -177 308 -173
rect 413 -171 418 -169
rect 422 -171 434 -169
rect 438 -171 442 -169
rect 446 -171 570 -169
rect 312 -176 343 -174
rect 363 -176 373 -174
rect 383 -176 385 -174
rect 265 -179 268 -177
rect 272 -179 290 -177
rect 294 -179 296 -177
rect 303 -178 309 -177
rect 199 -186 201 -182
rect 212 -188 214 -179
rect 220 -187 222 -185
rect 226 -187 236 -185
rect 240 -187 243 -185
rect 191 -210 193 -198
rect 191 -234 193 -214
rect 199 -218 201 -190
rect 303 -181 309 -180
rect 413 -179 458 -177
rect 462 -179 570 -177
rect 303 -185 308 -181
rect 312 -184 313 -182
rect 333 -184 393 -182
rect 403 -184 405 -182
rect 247 -187 276 -185
rect 280 -187 290 -185
rect 294 -187 296 -185
rect 303 -186 309 -185
rect 212 -195 222 -193
rect 226 -195 247 -193
rect 251 -195 253 -193
rect 303 -189 309 -188
rect 303 -193 308 -189
rect 413 -187 482 -185
rect 486 -187 538 -185
rect 542 -187 570 -185
rect 312 -192 343 -190
rect 363 -192 373 -190
rect 383 -192 385 -190
rect 265 -195 268 -193
rect 272 -195 290 -193
rect 294 -195 296 -193
rect 303 -194 309 -193
rect 212 -204 214 -195
rect 220 -203 222 -201
rect 226 -203 236 -201
rect 240 -203 243 -201
rect 303 -197 309 -196
rect 413 -195 506 -193
rect 510 -195 538 -193
rect 542 -195 570 -193
rect 303 -201 308 -197
rect 312 -200 313 -198
rect 333 -200 393 -198
rect 403 -200 405 -198
rect 247 -203 276 -201
rect 280 -203 290 -201
rect 294 -203 296 -201
rect 303 -202 309 -201
rect 212 -211 222 -209
rect 226 -211 247 -209
rect 251 -211 253 -209
rect 303 -205 309 -204
rect 303 -209 308 -205
rect 413 -203 450 -201
rect 454 -203 570 -201
rect 312 -208 343 -206
rect 363 -208 373 -206
rect 383 -208 385 -206
rect 265 -211 268 -209
rect 272 -211 290 -209
rect 294 -211 296 -209
rect 303 -210 309 -209
rect 212 -220 214 -211
rect 220 -219 222 -217
rect 226 -219 236 -217
rect 240 -219 243 -217
rect 183 -258 185 -238
rect 191 -258 193 -238
rect 167 -274 169 -270
rect 175 -274 177 -270
rect 151 -314 153 -310
rect 159 -314 161 -286
rect 167 -290 169 -278
rect 175 -290 177 -278
rect 183 -282 185 -262
rect 191 -282 193 -262
rect 199 -266 201 -222
rect 303 -213 309 -212
rect 413 -211 458 -209
rect 462 -211 570 -209
rect 303 -217 308 -213
rect 312 -216 313 -214
rect 333 -216 393 -214
rect 403 -216 405 -214
rect 247 -219 276 -217
rect 280 -219 290 -217
rect 294 -219 296 -217
rect 303 -218 309 -217
rect 212 -227 222 -225
rect 226 -227 247 -225
rect 251 -227 253 -225
rect 303 -221 309 -220
rect 303 -225 308 -221
rect 413 -219 426 -217
rect 430 -219 570 -217
rect 312 -224 343 -222
rect 363 -224 373 -222
rect 383 -224 385 -222
rect 265 -227 268 -225
rect 272 -227 290 -225
rect 294 -227 296 -225
rect 303 -226 309 -225
rect 212 -236 214 -227
rect 303 -229 309 -228
rect 413 -227 442 -225
rect 446 -227 570 -225
rect 303 -233 308 -229
rect 312 -232 313 -230
rect 333 -232 393 -230
rect 403 -232 405 -230
rect 303 -234 309 -233
rect 413 -235 482 -233
rect 486 -235 538 -233
rect 542 -235 570 -233
rect 220 -251 222 -249
rect 226 -251 236 -249
rect 240 -251 243 -249
rect 247 -251 276 -249
rect 280 -251 290 -249
rect 294 -251 296 -249
rect 212 -259 222 -257
rect 226 -259 247 -257
rect 251 -259 253 -257
rect 303 -253 309 -252
rect 303 -257 308 -253
rect 312 -256 343 -254
rect 363 -256 373 -254
rect 383 -256 385 -254
rect 265 -259 268 -257
rect 272 -259 290 -257
rect 294 -259 296 -257
rect 303 -258 309 -257
rect 212 -268 214 -259
rect 220 -267 222 -265
rect 226 -267 236 -265
rect 240 -267 243 -265
rect 199 -274 201 -270
rect 303 -261 309 -260
rect 413 -259 426 -257
rect 430 -259 570 -257
rect 303 -265 308 -261
rect 312 -264 313 -262
rect 333 -264 393 -262
rect 403 -264 405 -262
rect 247 -267 276 -265
rect 280 -267 290 -265
rect 294 -267 296 -265
rect 303 -266 309 -265
rect 212 -275 222 -273
rect 226 -275 247 -273
rect 251 -275 253 -273
rect 303 -269 309 -268
rect 303 -273 308 -269
rect 413 -267 506 -265
rect 510 -267 538 -265
rect 542 -267 570 -265
rect 312 -272 343 -270
rect 363 -272 373 -270
rect 383 -272 385 -270
rect 265 -275 268 -273
rect 272 -275 290 -273
rect 294 -275 296 -273
rect 303 -274 309 -273
rect 167 -306 169 -294
rect 135 -330 137 -326
rect 135 -338 137 -334
rect 143 -338 145 -326
rect 135 -346 137 -342
rect 135 -354 137 -350
rect 143 -354 145 -342
rect 135 -368 137 -358
rect 143 -368 145 -358
rect 151 -368 153 -318
rect 159 -330 161 -318
rect 159 -368 161 -334
rect 167 -338 169 -310
rect 167 -368 169 -342
rect 175 -346 177 -294
rect 183 -298 185 -286
rect 191 -290 193 -286
rect 183 -306 185 -302
rect 183 -322 185 -310
rect 191 -314 193 -294
rect 199 -298 201 -278
rect 212 -284 214 -275
rect 220 -283 222 -281
rect 226 -283 236 -281
rect 240 -283 243 -281
rect 303 -277 309 -276
rect 413 -275 426 -273
rect 430 -275 570 -273
rect 303 -281 308 -277
rect 312 -280 313 -278
rect 333 -280 393 -278
rect 403 -280 405 -278
rect 247 -283 276 -281
rect 280 -283 290 -281
rect 294 -283 296 -281
rect 303 -282 309 -281
rect 212 -291 222 -289
rect 226 -291 247 -289
rect 251 -291 253 -289
rect 303 -285 309 -284
rect 303 -289 308 -285
rect 413 -283 426 -281
rect 430 -283 434 -281
rect 438 -283 570 -281
rect 312 -288 343 -286
rect 363 -288 373 -286
rect 383 -288 385 -286
rect 265 -291 268 -289
rect 272 -291 290 -289
rect 294 -291 296 -289
rect 303 -290 309 -289
rect 212 -300 214 -291
rect 220 -299 222 -297
rect 226 -299 236 -297
rect 240 -299 243 -297
rect 175 -368 177 -350
rect 183 -368 185 -326
rect 191 -368 193 -318
rect 199 -330 201 -302
rect 303 -293 309 -292
rect 413 -291 434 -289
rect 438 -291 570 -289
rect 303 -297 308 -293
rect 312 -296 313 -294
rect 333 -296 393 -294
rect 403 -296 405 -294
rect 247 -299 276 -297
rect 280 -299 290 -297
rect 294 -299 296 -297
rect 303 -298 309 -297
rect 212 -307 222 -305
rect 226 -307 247 -305
rect 251 -307 253 -305
rect 303 -301 309 -300
rect 303 -305 308 -301
rect 413 -299 458 -297
rect 462 -299 570 -297
rect 312 -304 343 -302
rect 363 -304 373 -302
rect 383 -304 385 -302
rect 265 -307 268 -305
rect 272 -307 290 -305
rect 294 -307 296 -305
rect 303 -306 309 -305
rect 212 -316 214 -307
rect 220 -315 222 -313
rect 226 -315 236 -313
rect 240 -315 243 -313
rect 303 -309 309 -308
rect 413 -307 546 -305
rect 550 -307 570 -305
rect 303 -313 308 -309
rect 312 -312 313 -310
rect 333 -312 393 -310
rect 403 -312 405 -310
rect 247 -315 276 -313
rect 280 -315 290 -313
rect 294 -315 296 -313
rect 303 -314 309 -313
rect 212 -323 222 -321
rect 226 -323 247 -321
rect 251 -323 253 -321
rect 303 -317 309 -316
rect 303 -321 308 -317
rect 413 -315 538 -313
rect 542 -315 554 -313
rect 558 -315 570 -313
rect 312 -320 343 -318
rect 363 -320 373 -318
rect 383 -320 385 -318
rect 265 -323 268 -321
rect 272 -323 290 -321
rect 294 -323 296 -321
rect 303 -322 309 -321
rect 212 -332 214 -323
rect 220 -331 222 -329
rect 226 -331 236 -329
rect 240 -331 243 -329
rect 199 -346 201 -334
rect 303 -325 309 -324
rect 413 -323 442 -321
rect 446 -323 570 -321
rect 303 -329 308 -325
rect 312 -328 313 -326
rect 333 -328 393 -326
rect 403 -328 405 -326
rect 247 -331 276 -329
rect 280 -331 290 -329
rect 294 -331 296 -329
rect 303 -330 309 -329
rect 212 -339 222 -337
rect 226 -339 247 -337
rect 251 -339 253 -337
rect 303 -333 309 -332
rect 303 -337 308 -333
rect 413 -331 434 -329
rect 438 -331 570 -329
rect 312 -336 343 -334
rect 363 -336 373 -334
rect 383 -336 385 -334
rect 265 -339 268 -337
rect 272 -339 290 -337
rect 294 -339 296 -337
rect 303 -338 309 -337
rect 212 -348 214 -339
rect 303 -341 309 -340
rect 413 -339 442 -337
rect 446 -339 570 -337
rect 303 -345 308 -341
rect 312 -344 313 -342
rect 333 -344 393 -342
rect 403 -344 405 -342
rect 247 -347 276 -345
rect 280 -347 290 -345
rect 294 -347 296 -345
rect 303 -346 309 -345
rect 199 -354 201 -350
rect 303 -349 309 -348
rect 303 -353 308 -349
rect 413 -347 418 -345
rect 422 -347 570 -345
rect 312 -352 343 -350
rect 363 -352 373 -350
rect 383 -352 385 -350
rect 265 -355 268 -353
rect 272 -355 290 -353
rect 294 -355 296 -353
rect 303 -354 309 -353
rect 199 -368 201 -358
rect 413 -355 418 -353
rect 422 -355 442 -353
rect 446 -355 570 -353
rect 430 -366 433 -364
rect 446 -366 449 -364
rect 462 -366 465 -364
rect 478 -366 481 -364
rect 494 -366 497 -364
rect 518 -366 521 -364
rect 534 -366 537 -364
rect 550 -366 553 -364
rect 31 -370 32 -368
rect 39 -370 40 -368
rect 47 -370 48 -368
rect 55 -370 56 -368
rect 63 -370 64 -368
rect 71 -370 72 -368
rect 79 -370 80 -368
rect 87 -370 88 -368
rect 95 -370 96 -368
rect 103 -370 104 -368
rect 111 -370 112 -368
rect 119 -370 120 -368
rect 127 -370 128 -368
rect 135 -370 136 -368
rect 143 -370 144 -368
rect 151 -370 152 -368
rect 159 -370 160 -368
rect 167 -370 168 -368
rect 175 -370 176 -368
rect 183 -370 184 -368
rect 191 -370 192 -368
rect 199 -370 200 -368
rect 431 -376 433 -366
rect 37 -378 39 -376
rect 53 -378 55 -376
rect 69 -378 71 -376
rect 85 -378 87 -376
rect 101 -378 103 -376
rect 117 -378 119 -376
rect 133 -378 135 -376
rect 149 -378 151 -376
rect 165 -378 167 -376
rect 181 -378 183 -376
rect 197 -378 199 -376
rect 29 -401 31 -399
rect 29 -425 31 -415
rect 29 -488 31 -451
rect 37 -461 39 -391
rect 45 -401 47 -399
rect 45 -425 47 -415
rect 37 -488 39 -487
rect 45 -488 47 -451
rect 53 -461 55 -391
rect 61 -401 63 -399
rect 61 -425 63 -415
rect 53 -488 55 -487
rect 61 -488 63 -451
rect 69 -461 71 -391
rect 77 -401 79 -399
rect 77 -425 79 -415
rect 69 -488 71 -487
rect 77 -488 79 -451
rect 85 -461 87 -391
rect 93 -401 95 -399
rect 93 -425 95 -415
rect 85 -488 87 -487
rect 93 -488 95 -451
rect 101 -461 103 -391
rect 109 -401 111 -399
rect 109 -425 111 -415
rect 101 -488 103 -487
rect 109 -488 111 -451
rect 117 -461 119 -391
rect 125 -401 127 -399
rect 125 -425 127 -415
rect 117 -488 119 -487
rect 125 -488 127 -451
rect 133 -461 135 -391
rect 141 -401 143 -399
rect 141 -425 143 -415
rect 133 -488 135 -487
rect 141 -488 143 -451
rect 149 -461 151 -391
rect 157 -401 159 -399
rect 157 -425 159 -415
rect 149 -488 151 -487
rect 157 -488 159 -451
rect 165 -461 167 -391
rect 173 -401 175 -399
rect 173 -425 175 -415
rect 165 -488 167 -487
rect 173 -488 175 -451
rect 181 -461 183 -391
rect 447 -376 449 -366
rect 423 -391 425 -390
rect 189 -401 191 -399
rect 189 -425 191 -415
rect 181 -488 183 -487
rect 189 -488 191 -451
rect 197 -461 199 -391
rect 423 -405 425 -403
rect 423 -413 425 -411
rect 423 -438 425 -437
rect 431 -440 433 -388
rect 463 -376 465 -366
rect 439 -391 441 -390
rect 439 -405 441 -403
rect 439 -413 441 -411
rect 439 -438 441 -437
rect 197 -488 199 -487
rect 29 -490 30 -488
rect 37 -491 38 -488
rect 45 -490 46 -488
rect 53 -491 54 -488
rect 61 -490 62 -488
rect 69 -491 70 -488
rect 77 -490 78 -488
rect 85 -491 86 -488
rect 93 -490 94 -488
rect 101 -491 102 -488
rect 109 -490 110 -488
rect 117 -491 118 -488
rect 125 -490 126 -488
rect 133 -491 134 -488
rect 141 -490 142 -488
rect 149 -491 150 -488
rect 157 -490 158 -488
rect 165 -491 166 -488
rect 173 -490 174 -488
rect 181 -491 182 -488
rect 189 -490 190 -488
rect 197 -491 198 -488
rect 35 -505 38 -503
rect 42 -505 44 -503
rect 51 -505 54 -503
rect 58 -505 60 -503
rect 67 -505 70 -503
rect 74 -505 76 -503
rect 83 -505 86 -503
rect 90 -505 92 -503
rect 99 -505 102 -503
rect 106 -505 108 -503
rect 115 -505 118 -503
rect 122 -505 124 -503
rect 131 -505 134 -503
rect 138 -505 140 -503
rect 147 -505 150 -503
rect 154 -505 156 -503
rect 163 -505 166 -503
rect 170 -505 172 -503
rect 179 -505 182 -503
rect 186 -505 188 -503
rect 195 -505 198 -503
rect 202 -505 204 -503
rect 35 -510 38 -508
rect 42 -510 44 -508
rect 51 -510 54 -508
rect 58 -510 60 -508
rect 67 -510 70 -508
rect 74 -510 76 -508
rect 83 -510 86 -508
rect 90 -510 92 -508
rect 99 -510 102 -508
rect 106 -510 108 -508
rect 115 -510 118 -508
rect 122 -510 124 -508
rect 131 -510 134 -508
rect 138 -510 140 -508
rect 147 -510 150 -508
rect 154 -510 156 -508
rect 163 -510 166 -508
rect 170 -510 172 -508
rect 179 -510 182 -508
rect 186 -510 188 -508
rect 195 -510 198 -508
rect 202 -510 204 -508
rect 423 -509 425 -442
rect 447 -440 449 -388
rect 479 -376 481 -366
rect 455 -391 457 -390
rect 455 -405 457 -403
rect 455 -413 457 -411
rect 455 -438 457 -437
rect 431 -466 433 -464
rect 431 -481 433 -478
rect 35 -518 37 -510
rect 51 -518 53 -510
rect 67 -518 69 -510
rect 83 -518 85 -510
rect 99 -518 101 -510
rect 115 -518 117 -510
rect 131 -518 133 -510
rect 147 -518 149 -510
rect 163 -518 165 -510
rect 179 -518 181 -510
rect 195 -518 197 -510
rect 35 -536 38 -534
rect 42 -536 44 -534
rect 51 -536 54 -534
rect 58 -536 60 -534
rect 67 -536 70 -534
rect 74 -536 76 -534
rect 83 -536 86 -534
rect 90 -536 92 -534
rect 99 -536 102 -534
rect 106 -536 108 -534
rect 115 -536 118 -534
rect 122 -536 124 -534
rect 131 -536 134 -534
rect 138 -536 140 -534
rect 147 -536 150 -534
rect 154 -536 156 -534
rect 163 -536 166 -534
rect 170 -536 172 -534
rect 179 -536 182 -534
rect 186 -536 188 -534
rect 195 -536 198 -534
rect 202 -536 204 -534
rect 423 -535 425 -533
rect 35 -541 38 -539
rect 42 -541 44 -539
rect 51 -541 54 -539
rect 58 -541 60 -539
rect 67 -541 70 -539
rect 74 -541 76 -539
rect 83 -541 86 -539
rect 90 -541 92 -539
rect 99 -541 102 -539
rect 106 -541 108 -539
rect 115 -541 118 -539
rect 122 -541 124 -539
rect 131 -541 134 -539
rect 138 -541 140 -539
rect 147 -541 150 -539
rect 154 -541 156 -539
rect 163 -541 166 -539
rect 170 -541 172 -539
rect 179 -541 182 -539
rect 186 -541 188 -539
rect 195 -541 198 -539
rect 202 -541 204 -539
rect 35 -549 37 -541
rect 51 -549 53 -541
rect 67 -549 69 -541
rect 83 -549 85 -541
rect 99 -549 101 -541
rect 115 -549 117 -541
rect 131 -549 133 -541
rect 147 -549 149 -541
rect 163 -549 165 -541
rect 179 -549 181 -541
rect 195 -549 197 -541
rect 423 -543 425 -541
rect 35 -561 37 -553
rect 51 -561 53 -553
rect 67 -561 69 -553
rect 83 -561 85 -553
rect 99 -561 101 -553
rect 115 -561 117 -553
rect 131 -561 133 -553
rect 147 -561 149 -553
rect 163 -561 165 -553
rect 179 -561 181 -553
rect 195 -561 197 -553
rect 423 -556 425 -555
rect 431 -558 433 -505
rect 439 -509 441 -442
rect 463 -440 465 -388
rect 495 -376 497 -366
rect 471 -391 473 -390
rect 471 -405 473 -403
rect 471 -413 473 -411
rect 471 -438 473 -437
rect 447 -466 449 -464
rect 447 -481 449 -478
rect 439 -535 441 -533
rect 439 -543 441 -541
rect 439 -556 441 -555
rect 35 -563 38 -561
rect 42 -563 44 -561
rect 51 -563 54 -561
rect 58 -563 60 -561
rect 67 -563 70 -561
rect 74 -563 76 -561
rect 83 -563 86 -561
rect 90 -563 92 -561
rect 99 -563 102 -561
rect 106 -563 108 -561
rect 115 -563 118 -561
rect 122 -563 124 -561
rect 131 -563 134 -561
rect 138 -563 140 -561
rect 147 -563 150 -561
rect 154 -563 156 -561
rect 163 -563 166 -561
rect 170 -563 172 -561
rect 179 -563 182 -561
rect 186 -563 188 -561
rect 195 -563 198 -561
rect 202 -563 204 -561
rect 35 -568 38 -566
rect 42 -568 44 -566
rect 51 -568 54 -566
rect 58 -568 60 -566
rect 67 -568 70 -566
rect 74 -568 76 -566
rect 83 -568 86 -566
rect 90 -568 92 -566
rect 99 -568 102 -566
rect 106 -568 108 -566
rect 115 -568 118 -566
rect 122 -568 124 -566
rect 131 -568 134 -566
rect 138 -568 140 -566
rect 147 -568 150 -566
rect 154 -568 156 -566
rect 163 -568 166 -566
rect 170 -568 172 -566
rect 179 -568 182 -566
rect 186 -568 188 -566
rect 195 -568 198 -566
rect 202 -568 204 -566
rect 447 -558 449 -505
rect 455 -509 457 -442
rect 479 -440 481 -388
rect 519 -376 521 -366
rect 487 -391 489 -390
rect 487 -405 489 -403
rect 487 -413 489 -411
rect 487 -438 489 -437
rect 463 -466 465 -464
rect 463 -481 465 -478
rect 455 -535 457 -533
rect 455 -543 457 -541
rect 455 -556 457 -555
rect 431 -572 433 -570
rect 463 -558 465 -505
rect 471 -509 473 -442
rect 495 -440 497 -388
rect 535 -376 537 -366
rect 511 -391 513 -390
rect 511 -405 513 -403
rect 511 -413 513 -411
rect 511 -438 513 -437
rect 479 -466 481 -464
rect 479 -481 481 -478
rect 471 -535 473 -533
rect 471 -543 473 -541
rect 471 -556 473 -555
rect 447 -572 449 -570
rect 479 -558 481 -505
rect 487 -509 489 -442
rect 519 -440 521 -388
rect 551 -376 553 -366
rect 527 -391 529 -390
rect 527 -405 529 -403
rect 527 -413 529 -411
rect 527 -438 529 -437
rect 495 -466 497 -464
rect 495 -481 497 -478
rect 487 -535 489 -533
rect 487 -543 489 -541
rect 487 -556 489 -555
rect 463 -572 465 -570
rect 495 -558 497 -505
rect 511 -509 513 -442
rect 535 -440 537 -388
rect 543 -391 545 -390
rect 543 -405 545 -403
rect 543 -413 545 -411
rect 543 -438 545 -437
rect 519 -466 521 -464
rect 519 -481 521 -478
rect 511 -535 513 -533
rect 511 -543 513 -541
rect 511 -556 513 -555
rect 479 -572 481 -570
rect 519 -558 521 -505
rect 527 -509 529 -442
rect 551 -440 553 -388
rect 535 -466 537 -464
rect 535 -481 537 -478
rect 527 -535 529 -533
rect 527 -543 529 -541
rect 527 -556 529 -555
rect 495 -572 497 -570
rect 535 -558 537 -505
rect 543 -509 545 -442
rect 551 -466 553 -464
rect 551 -481 553 -478
rect 543 -535 545 -533
rect 543 -543 545 -541
rect 543 -556 545 -555
rect 519 -572 521 -570
rect 551 -558 553 -505
rect 559 -509 561 -442
rect 567 -481 569 -478
rect 559 -535 561 -533
rect 559 -543 561 -541
rect 559 -556 561 -555
rect 535 -572 537 -570
rect 567 -558 569 -505
rect 551 -572 553 -570
rect 567 -572 569 -570
<< ndiffusion >>
rect 34 -2 38 1
rect 34 -6 39 -2
rect 41 -6 42 -2
rect 34 -10 38 -6
rect 34 -14 39 -10
rect 41 -14 42 -10
rect 34 -18 38 -14
rect 50 -10 54 1
rect 66 -10 70 1
rect 50 -14 55 -10
rect 57 -14 58 -10
rect 62 -14 63 -10
rect 65 -14 70 -10
rect 50 -18 54 -14
rect 34 -22 39 -18
rect 41 -22 42 -18
rect 46 -22 47 -18
rect 49 -22 54 -18
rect 34 -26 38 -22
rect 34 -30 39 -26
rect 41 -30 42 -26
rect 34 -34 38 -30
rect 34 -38 39 -34
rect 41 -38 42 -34
rect 34 -42 38 -38
rect 34 -46 39 -42
rect 41 -46 42 -42
rect 34 -50 38 -46
rect 34 -54 39 -50
rect 41 -54 42 -50
rect 34 -58 38 -54
rect 34 -62 39 -58
rect 41 -62 42 -58
rect 34 -66 38 -62
rect 34 -70 39 -66
rect 41 -70 42 -66
rect 34 -74 38 -70
rect 34 -78 39 -74
rect 41 -78 42 -74
rect 34 -82 38 -78
rect 34 -86 39 -82
rect 41 -86 42 -82
rect 34 -114 38 -86
rect 34 -154 38 -118
rect 34 -158 39 -154
rect 41 -158 42 -154
rect 34 -162 38 -158
rect 50 -34 54 -22
rect 50 -38 55 -34
rect 57 -38 58 -34
rect 50 -114 54 -38
rect 50 -162 54 -118
rect 34 -166 39 -162
rect 41 -166 42 -162
rect 46 -166 47 -162
rect 49 -166 54 -162
rect 34 -170 38 -166
rect 34 -174 39 -170
rect 41 -174 42 -170
rect 34 -202 38 -174
rect 34 -206 39 -202
rect 41 -206 42 -202
rect 34 -218 38 -206
rect 34 -222 39 -218
rect 41 -222 42 -218
rect 34 -226 38 -222
rect 34 -230 39 -226
rect 41 -230 42 -226
rect 34 -242 38 -230
rect 34 -258 38 -246
rect 34 -262 39 -258
rect 41 -262 42 -258
rect 34 -274 38 -262
rect 34 -278 39 -274
rect 41 -278 42 -274
rect 34 -282 38 -278
rect 34 -286 39 -282
rect 41 -286 42 -282
rect 34 -290 38 -286
rect 34 -294 39 -290
rect 41 -294 42 -290
rect 34 -322 38 -294
rect 34 -326 39 -322
rect 41 -326 42 -322
rect 34 -330 38 -326
rect 34 -334 39 -330
rect 41 -334 42 -330
rect 34 -338 38 -334
rect 34 -342 39 -338
rect 41 -342 42 -338
rect 34 -346 38 -342
rect 34 -350 39 -346
rect 41 -350 42 -346
rect 34 -354 38 -350
rect 34 -358 39 -354
rect 41 -358 42 -354
rect 34 -361 38 -358
rect 50 -242 54 -166
rect 50 -361 54 -246
rect 66 -18 70 -14
rect 66 -22 71 -18
rect 73 -22 74 -18
rect 66 -114 70 -22
rect 66 -154 70 -118
rect 62 -158 63 -154
rect 65 -158 70 -154
rect 66 -242 70 -158
rect 66 -361 70 -246
rect 82 -26 86 1
rect 78 -30 79 -26
rect 81 -30 86 -26
rect 82 -58 86 -30
rect 98 -2 102 1
rect 114 -2 118 1
rect 98 -6 103 -2
rect 105 -6 106 -2
rect 110 -6 111 -2
rect 113 -6 118 -2
rect 98 -50 102 -6
rect 94 -54 95 -50
rect 97 -54 102 -50
rect 82 -62 87 -58
rect 89 -62 90 -58
rect 82 -74 86 -62
rect 82 -78 87 -74
rect 89 -78 90 -74
rect 82 -114 86 -78
rect 82 -242 86 -118
rect 82 -361 86 -246
rect 98 -114 102 -54
rect 98 -242 102 -118
rect 98 -361 102 -246
rect 114 -42 118 -6
rect 130 -2 134 1
rect 126 -6 127 -2
rect 129 -6 134 -2
rect 130 -10 134 -6
rect 130 -14 135 -10
rect 137 -14 138 -10
rect 130 -18 134 -14
rect 130 -22 135 -18
rect 137 -22 138 -18
rect 130 -34 134 -22
rect 146 -2 150 1
rect 146 -6 151 -2
rect 153 -6 154 -2
rect 146 -10 150 -6
rect 146 -14 151 -10
rect 153 -14 154 -10
rect 146 -26 150 -14
rect 146 -30 151 -26
rect 153 -30 154 -26
rect 146 -34 150 -30
rect 130 -38 135 -34
rect 137 -38 138 -34
rect 142 -38 143 -34
rect 145 -38 150 -34
rect 130 -42 134 -38
rect 114 -46 119 -42
rect 121 -46 122 -42
rect 126 -46 127 -42
rect 129 -46 134 -42
rect 114 -114 118 -46
rect 114 -242 118 -118
rect 114 -361 118 -246
rect 130 -50 134 -46
rect 126 -54 127 -50
rect 129 -54 134 -50
rect 130 -58 134 -54
rect 126 -62 127 -58
rect 129 -62 134 -58
rect 130 -66 134 -62
rect 146 -42 150 -38
rect 146 -46 151 -42
rect 153 -46 154 -42
rect 146 -50 150 -46
rect 146 -54 151 -50
rect 153 -54 154 -50
rect 146 -58 150 -54
rect 162 -2 166 1
rect 162 -6 167 -2
rect 169 -6 170 -2
rect 162 -10 166 -6
rect 162 -14 167 -10
rect 169 -14 170 -10
rect 162 -18 166 -14
rect 162 -22 167 -18
rect 169 -22 170 -18
rect 162 -26 166 -22
rect 178 -2 182 1
rect 178 -6 183 -2
rect 185 -6 186 -2
rect 178 -10 182 -6
rect 178 -14 183 -10
rect 185 -14 186 -10
rect 178 -26 182 -14
rect 162 -30 167 -26
rect 169 -30 170 -26
rect 174 -30 175 -26
rect 177 -30 182 -26
rect 162 -34 166 -30
rect 162 -38 167 -34
rect 169 -38 170 -34
rect 162 -42 166 -38
rect 162 -46 167 -42
rect 169 -46 170 -42
rect 162 -50 166 -46
rect 162 -54 167 -50
rect 169 -54 170 -50
rect 162 -58 166 -54
rect 146 -62 151 -58
rect 153 -62 154 -58
rect 158 -62 159 -58
rect 161 -62 166 -58
rect 146 -66 150 -62
rect 130 -70 135 -66
rect 137 -70 138 -66
rect 142 -70 143 -66
rect 145 -70 150 -66
rect 130 -74 134 -70
rect 126 -78 127 -74
rect 129 -78 134 -74
rect 130 -82 134 -78
rect 126 -86 127 -82
rect 129 -86 134 -82
rect 130 -90 134 -86
rect 126 -94 127 -90
rect 129 -94 134 -90
rect 130 -98 134 -94
rect 146 -74 150 -70
rect 162 -66 166 -62
rect 158 -70 159 -66
rect 161 -70 166 -66
rect 146 -78 151 -74
rect 153 -78 154 -74
rect 146 -82 150 -78
rect 162 -74 166 -70
rect 178 -34 182 -30
rect 194 -2 198 1
rect 236 7 240 8
rect 236 3 240 5
rect 276 7 280 8
rect 276 3 280 5
rect 236 0 251 3
rect 247 -1 251 0
rect 194 -6 199 -2
rect 201 -6 202 -2
rect 268 0 280 3
rect 268 -1 272 0
rect 373 2 383 3
rect 194 -10 198 -6
rect 194 -14 199 -10
rect 201 -14 202 -10
rect 247 -4 251 -3
rect 268 -4 272 -3
rect 247 -7 250 -4
rect 236 -9 240 -8
rect 194 -18 198 -14
rect 236 -13 240 -11
rect 276 -9 280 -8
rect 373 -1 383 0
rect 418 -1 422 0
rect 450 -1 454 0
rect 401 -5 403 -1
rect 418 -4 422 -3
rect 450 -4 454 -3
rect 393 -6 403 -5
rect 414 -8 498 -4
rect 502 -8 563 -4
rect 393 -9 403 -8
rect 418 -9 422 -8
rect 426 -9 430 -8
rect 434 -9 438 -8
rect 276 -13 280 -11
rect 236 -16 251 -13
rect 247 -17 251 -16
rect 194 -22 199 -18
rect 201 -22 202 -18
rect 268 -16 280 -13
rect 268 -17 272 -16
rect 418 -12 422 -11
rect 373 -14 383 -13
rect 426 -12 430 -11
rect 434 -12 438 -11
rect 194 -26 198 -22
rect 190 -30 191 -26
rect 193 -30 198 -26
rect 178 -38 183 -34
rect 185 -38 186 -34
rect 178 -58 182 -38
rect 178 -62 183 -58
rect 185 -62 186 -58
rect 178 -66 182 -62
rect 174 -70 175 -66
rect 177 -70 182 -66
rect 178 -74 182 -70
rect 162 -78 167 -74
rect 169 -78 170 -74
rect 174 -78 175 -74
rect 177 -78 182 -74
rect 162 -82 166 -78
rect 146 -86 151 -82
rect 153 -86 154 -82
rect 158 -86 159 -82
rect 161 -86 166 -82
rect 146 -90 150 -86
rect 162 -90 166 -86
rect 146 -94 151 -90
rect 153 -94 154 -90
rect 158 -94 159 -90
rect 161 -94 166 -90
rect 146 -98 150 -94
rect 130 -102 135 -98
rect 137 -102 138 -98
rect 142 -102 143 -98
rect 145 -102 150 -98
rect 130 -106 134 -102
rect 146 -106 150 -102
rect 130 -110 135 -106
rect 137 -110 138 -106
rect 142 -110 143 -106
rect 145 -110 150 -106
rect 130 -114 134 -110
rect 130 -130 134 -118
rect 146 -114 150 -110
rect 146 -130 150 -118
rect 130 -134 135 -130
rect 137 -134 138 -130
rect 142 -134 143 -130
rect 145 -134 150 -130
rect 130 -138 134 -134
rect 126 -142 127 -138
rect 129 -142 134 -138
rect 130 -146 134 -142
rect 126 -150 127 -146
rect 129 -150 134 -146
rect 130 -154 134 -150
rect 130 -158 135 -154
rect 137 -158 138 -154
rect 130 -162 134 -158
rect 130 -166 135 -162
rect 137 -166 138 -162
rect 130 -170 134 -166
rect 126 -174 127 -170
rect 129 -174 134 -170
rect 130 -178 134 -174
rect 130 -182 135 -178
rect 137 -182 138 -178
rect 130 -186 134 -182
rect 146 -138 150 -134
rect 162 -98 166 -94
rect 158 -102 159 -98
rect 161 -102 166 -98
rect 162 -106 166 -102
rect 158 -110 159 -106
rect 161 -110 166 -106
rect 162 -114 166 -110
rect 162 -130 166 -118
rect 158 -134 159 -130
rect 161 -134 166 -130
rect 146 -142 151 -138
rect 153 -142 154 -138
rect 146 -146 150 -142
rect 146 -150 151 -146
rect 153 -150 154 -146
rect 146 -170 150 -150
rect 162 -138 166 -134
rect 178 -82 182 -78
rect 194 -42 198 -30
rect 247 -20 251 -19
rect 268 -20 272 -19
rect 247 -23 250 -20
rect 236 -25 240 -24
rect 236 -29 240 -27
rect 276 -25 280 -24
rect 373 -17 383 -16
rect 418 -17 422 -16
rect 401 -21 403 -17
rect 418 -20 422 -19
rect 393 -22 403 -21
rect 414 -24 498 -20
rect 502 -24 563 -20
rect 393 -25 403 -24
rect 434 -25 438 -24
rect 276 -29 280 -27
rect 236 -32 251 -29
rect 247 -33 251 -32
rect 268 -32 280 -29
rect 268 -33 272 -32
rect 434 -28 438 -27
rect 373 -30 383 -29
rect 194 -46 199 -42
rect 201 -46 202 -42
rect 247 -36 251 -35
rect 268 -36 272 -35
rect 247 -39 250 -36
rect 236 -41 240 -40
rect 194 -50 198 -46
rect 236 -45 240 -43
rect 276 -41 280 -40
rect 373 -33 383 -32
rect 418 -33 422 -32
rect 401 -37 403 -33
rect 418 -36 422 -35
rect 393 -38 403 -37
rect 414 -40 498 -36
rect 502 -40 563 -36
rect 393 -41 403 -40
rect 426 -41 430 -40
rect 450 -41 454 -40
rect 276 -45 280 -43
rect 236 -48 251 -45
rect 247 -49 251 -48
rect 194 -54 199 -50
rect 201 -54 202 -50
rect 268 -48 280 -45
rect 268 -49 272 -48
rect 426 -44 430 -43
rect 373 -46 383 -45
rect 194 -66 198 -54
rect 190 -70 191 -66
rect 193 -70 198 -66
rect 178 -86 183 -82
rect 185 -86 186 -82
rect 178 -90 182 -86
rect 194 -82 198 -70
rect 247 -52 251 -51
rect 268 -52 272 -51
rect 247 -55 250 -52
rect 236 -57 240 -56
rect 236 -61 240 -59
rect 276 -57 280 -56
rect 373 -49 383 -48
rect 426 -49 430 -48
rect 450 -44 454 -43
rect 450 -49 454 -48
rect 401 -53 403 -49
rect 426 -52 430 -51
rect 450 -52 454 -51
rect 393 -54 403 -53
rect 414 -56 498 -52
rect 502 -56 563 -52
rect 393 -57 403 -56
rect 418 -57 422 -56
rect 434 -57 438 -56
rect 450 -57 454 -56
rect 276 -61 280 -59
rect 236 -64 251 -61
rect 247 -65 251 -64
rect 268 -64 280 -61
rect 268 -65 272 -64
rect 418 -60 422 -59
rect 373 -62 383 -61
rect 434 -60 438 -59
rect 450 -60 454 -59
rect 247 -68 251 -67
rect 268 -68 272 -67
rect 247 -71 250 -68
rect 236 -73 240 -72
rect 236 -77 240 -75
rect 276 -73 280 -72
rect 373 -65 383 -64
rect 450 -65 454 -64
rect 401 -69 403 -65
rect 450 -68 454 -67
rect 393 -70 403 -69
rect 414 -72 498 -68
rect 502 -72 563 -68
rect 393 -73 403 -72
rect 418 -73 422 -72
rect 426 -73 430 -72
rect 276 -77 280 -75
rect 236 -80 251 -77
rect 247 -81 251 -80
rect 194 -86 199 -82
rect 201 -86 202 -82
rect 268 -80 280 -77
rect 268 -81 272 -80
rect 418 -76 422 -75
rect 373 -78 383 -77
rect 426 -76 430 -75
rect 194 -90 198 -86
rect 178 -94 183 -90
rect 185 -94 186 -90
rect 190 -94 191 -90
rect 193 -94 198 -90
rect 178 -98 182 -94
rect 194 -98 198 -94
rect 178 -102 183 -98
rect 185 -102 186 -98
rect 190 -102 191 -98
rect 193 -102 198 -98
rect 178 -106 182 -102
rect 174 -110 175 -106
rect 177 -110 182 -106
rect 178 -114 182 -110
rect 178 -130 182 -118
rect 174 -134 175 -130
rect 177 -134 182 -130
rect 178 -138 182 -134
rect 162 -142 167 -138
rect 169 -142 170 -138
rect 174 -142 175 -138
rect 177 -142 182 -138
rect 162 -146 166 -142
rect 162 -150 167 -146
rect 169 -150 170 -146
rect 162 -154 166 -150
rect 158 -158 159 -154
rect 161 -158 166 -154
rect 146 -174 151 -170
rect 153 -174 154 -170
rect 146 -178 150 -174
rect 162 -170 166 -158
rect 162 -174 167 -170
rect 169 -174 170 -170
rect 162 -178 166 -174
rect 146 -182 151 -178
rect 153 -182 154 -178
rect 158 -182 159 -178
rect 161 -182 166 -178
rect 146 -186 150 -182
rect 130 -190 135 -186
rect 137 -190 138 -186
rect 142 -190 143 -186
rect 145 -190 150 -186
rect 130 -194 134 -190
rect 146 -194 150 -190
rect 130 -198 135 -194
rect 137 -198 138 -194
rect 142 -198 143 -194
rect 145 -198 150 -194
rect 130 -202 134 -198
rect 126 -206 127 -202
rect 129 -206 134 -202
rect 130 -210 134 -206
rect 130 -214 135 -210
rect 137 -214 138 -210
rect 130 -218 134 -214
rect 146 -202 150 -198
rect 146 -206 151 -202
rect 153 -206 154 -202
rect 146 -210 150 -206
rect 146 -214 151 -210
rect 153 -214 154 -210
rect 146 -218 150 -214
rect 130 -222 135 -218
rect 137 -222 138 -218
rect 142 -222 143 -218
rect 145 -222 150 -218
rect 130 -226 134 -222
rect 130 -230 135 -226
rect 137 -230 138 -226
rect 130 -234 134 -230
rect 130 -238 135 -234
rect 137 -238 138 -234
rect 130 -242 134 -238
rect 130 -266 134 -246
rect 130 -270 135 -266
rect 137 -270 138 -266
rect 130 -282 134 -270
rect 130 -286 135 -282
rect 137 -286 138 -282
rect 130 -290 134 -286
rect 130 -294 135 -290
rect 137 -294 138 -290
rect 130 -298 134 -294
rect 146 -226 150 -222
rect 162 -186 166 -182
rect 178 -146 182 -142
rect 194 -106 198 -102
rect 190 -110 191 -106
rect 193 -110 198 -106
rect 194 -114 198 -110
rect 194 -130 198 -118
rect 247 -84 251 -83
rect 268 -84 272 -83
rect 247 -87 250 -84
rect 236 -89 240 -88
rect 236 -93 240 -91
rect 276 -89 280 -88
rect 373 -81 383 -80
rect 434 -81 438 -80
rect 450 -81 454 -80
rect 401 -85 403 -81
rect 434 -84 438 -83
rect 450 -84 454 -83
rect 393 -86 403 -85
rect 414 -88 498 -84
rect 502 -88 563 -84
rect 393 -89 403 -88
rect 474 -89 478 -88
rect 490 -89 494 -88
rect 276 -93 280 -91
rect 236 -96 251 -93
rect 247 -97 251 -96
rect 268 -96 280 -93
rect 268 -97 272 -96
rect 474 -92 478 -91
rect 373 -94 383 -93
rect 490 -92 494 -91
rect 247 -100 251 -99
rect 268 -100 272 -99
rect 247 -103 250 -100
rect 373 -97 383 -96
rect 514 -97 518 -96
rect 401 -101 403 -97
rect 514 -100 518 -99
rect 393 -102 403 -101
rect 414 -104 498 -100
rect 502 -104 563 -100
rect 393 -105 403 -104
rect 546 -105 550 -104
rect 546 -108 550 -107
rect 236 -121 240 -120
rect 236 -125 240 -123
rect 276 -121 280 -120
rect 276 -125 280 -123
rect 236 -128 251 -125
rect 247 -129 251 -128
rect 194 -134 199 -130
rect 201 -134 202 -130
rect 268 -128 280 -125
rect 268 -129 272 -128
rect 373 -126 383 -125
rect 194 -138 198 -134
rect 190 -142 191 -138
rect 193 -142 198 -138
rect 194 -146 198 -142
rect 178 -150 183 -146
rect 185 -150 186 -146
rect 190 -150 191 -146
rect 193 -150 198 -146
rect 178 -162 182 -150
rect 194 -154 198 -150
rect 247 -132 251 -131
rect 268 -132 272 -131
rect 247 -135 250 -132
rect 236 -137 240 -136
rect 236 -141 240 -139
rect 276 -137 280 -136
rect 373 -129 383 -128
rect 530 -129 534 -128
rect 401 -133 403 -129
rect 530 -132 534 -131
rect 393 -134 403 -133
rect 414 -136 498 -132
rect 502 -136 563 -132
rect 393 -137 403 -136
rect 466 -137 470 -136
rect 522 -137 526 -136
rect 276 -141 280 -139
rect 236 -144 251 -141
rect 247 -145 251 -144
rect 268 -144 280 -141
rect 268 -145 272 -144
rect 466 -140 470 -139
rect 522 -140 526 -139
rect 373 -142 383 -141
rect 194 -158 199 -154
rect 201 -158 202 -154
rect 247 -148 251 -147
rect 268 -148 272 -147
rect 247 -151 250 -148
rect 236 -153 240 -152
rect 194 -162 198 -158
rect 178 -166 183 -162
rect 185 -166 186 -162
rect 190 -166 191 -162
rect 193 -166 198 -162
rect 178 -170 182 -166
rect 194 -170 198 -166
rect 178 -174 183 -170
rect 185 -174 186 -170
rect 190 -174 191 -170
rect 193 -174 198 -170
rect 178 -178 182 -174
rect 174 -182 175 -178
rect 177 -182 182 -178
rect 178 -186 182 -182
rect 162 -190 167 -186
rect 169 -190 170 -186
rect 174 -190 175 -186
rect 177 -190 182 -186
rect 162 -194 166 -190
rect 178 -194 182 -190
rect 162 -198 167 -194
rect 169 -198 170 -194
rect 174 -198 175 -194
rect 177 -198 182 -194
rect 162 -202 166 -198
rect 178 -202 182 -198
rect 162 -206 167 -202
rect 169 -206 170 -202
rect 174 -206 175 -202
rect 177 -206 182 -202
rect 162 -210 166 -206
rect 178 -210 182 -206
rect 162 -214 167 -210
rect 169 -214 170 -210
rect 174 -214 175 -210
rect 177 -214 182 -210
rect 162 -226 166 -214
rect 146 -230 151 -226
rect 153 -230 154 -226
rect 158 -230 159 -226
rect 161 -230 166 -226
rect 146 -234 150 -230
rect 146 -238 151 -234
rect 153 -238 154 -234
rect 146 -242 150 -238
rect 146 -258 150 -246
rect 146 -262 151 -258
rect 153 -262 154 -258
rect 146 -266 150 -262
rect 146 -270 151 -266
rect 153 -270 154 -266
rect 146 -274 150 -270
rect 146 -278 151 -274
rect 153 -278 154 -274
rect 146 -298 150 -278
rect 130 -302 135 -298
rect 137 -302 138 -298
rect 142 -302 143 -298
rect 145 -302 150 -298
rect 130 -306 134 -302
rect 126 -310 127 -306
rect 129 -310 134 -306
rect 130 -314 134 -310
rect 130 -318 135 -314
rect 137 -318 138 -314
rect 130 -322 134 -318
rect 146 -306 150 -302
rect 162 -234 166 -230
rect 178 -218 182 -214
rect 174 -222 175 -218
rect 177 -222 182 -218
rect 178 -226 182 -222
rect 174 -230 175 -226
rect 177 -230 182 -226
rect 162 -238 167 -234
rect 169 -238 170 -234
rect 162 -242 166 -238
rect 162 -258 166 -246
rect 162 -262 167 -258
rect 169 -262 170 -258
rect 162 -266 166 -262
rect 178 -234 182 -230
rect 194 -178 198 -174
rect 236 -157 240 -155
rect 276 -153 280 -152
rect 373 -145 383 -144
rect 506 -145 510 -144
rect 530 -145 534 -144
rect 401 -149 403 -145
rect 506 -148 510 -147
rect 530 -148 534 -147
rect 393 -150 403 -149
rect 414 -152 498 -148
rect 502 -152 563 -148
rect 393 -153 403 -152
rect 418 -153 422 -152
rect 276 -157 280 -155
rect 236 -160 251 -157
rect 247 -161 251 -160
rect 268 -160 280 -157
rect 268 -161 272 -160
rect 418 -156 422 -155
rect 373 -158 383 -157
rect 247 -164 251 -163
rect 268 -164 272 -163
rect 247 -167 250 -164
rect 236 -169 240 -168
rect 236 -173 240 -171
rect 276 -169 280 -168
rect 373 -161 383 -160
rect 426 -161 430 -160
rect 401 -165 403 -161
rect 426 -164 430 -163
rect 393 -166 403 -165
rect 414 -168 498 -164
rect 502 -168 563 -164
rect 393 -169 403 -168
rect 418 -169 422 -168
rect 434 -169 438 -168
rect 442 -169 446 -168
rect 276 -173 280 -171
rect 236 -176 251 -173
rect 247 -177 251 -176
rect 194 -182 199 -178
rect 201 -182 202 -178
rect 268 -176 280 -173
rect 268 -177 272 -176
rect 418 -172 422 -171
rect 373 -174 383 -173
rect 434 -172 438 -171
rect 442 -172 446 -171
rect 194 -186 198 -182
rect 194 -190 199 -186
rect 201 -190 202 -186
rect 247 -180 251 -179
rect 268 -180 272 -179
rect 247 -183 250 -180
rect 236 -185 240 -184
rect 194 -194 198 -190
rect 190 -198 191 -194
rect 193 -198 198 -194
rect 194 -210 198 -198
rect 190 -214 191 -210
rect 193 -214 198 -210
rect 194 -218 198 -214
rect 236 -189 240 -187
rect 276 -185 280 -184
rect 373 -177 383 -176
rect 458 -177 462 -176
rect 401 -181 403 -177
rect 458 -180 462 -179
rect 393 -182 403 -181
rect 414 -184 498 -180
rect 502 -184 563 -180
rect 393 -185 403 -184
rect 482 -185 486 -184
rect 538 -185 542 -184
rect 276 -189 280 -187
rect 236 -192 251 -189
rect 247 -193 251 -192
rect 268 -192 280 -189
rect 268 -193 272 -192
rect 482 -188 486 -187
rect 538 -188 542 -187
rect 373 -190 383 -189
rect 247 -196 251 -195
rect 268 -196 272 -195
rect 247 -199 250 -196
rect 236 -201 240 -200
rect 236 -205 240 -203
rect 276 -201 280 -200
rect 373 -193 383 -192
rect 506 -193 510 -192
rect 538 -193 542 -192
rect 401 -197 403 -193
rect 506 -196 510 -195
rect 538 -196 542 -195
rect 393 -198 403 -197
rect 414 -200 498 -196
rect 502 -200 563 -196
rect 393 -201 403 -200
rect 450 -201 454 -200
rect 276 -205 280 -203
rect 236 -208 251 -205
rect 247 -209 251 -208
rect 268 -208 280 -205
rect 268 -209 272 -208
rect 450 -204 454 -203
rect 373 -206 383 -205
rect 194 -222 199 -218
rect 201 -222 202 -218
rect 247 -212 251 -211
rect 268 -212 272 -211
rect 247 -215 250 -212
rect 236 -217 240 -216
rect 194 -234 198 -222
rect 178 -238 183 -234
rect 185 -238 186 -234
rect 190 -238 191 -234
rect 193 -238 198 -234
rect 178 -242 182 -238
rect 178 -258 182 -246
rect 194 -242 198 -238
rect 194 -258 198 -246
rect 178 -262 183 -258
rect 185 -262 186 -258
rect 190 -262 191 -258
rect 193 -262 198 -258
rect 178 -266 182 -262
rect 162 -270 167 -266
rect 169 -270 170 -266
rect 174 -270 175 -266
rect 177 -270 182 -266
rect 162 -274 166 -270
rect 178 -274 182 -270
rect 162 -278 167 -274
rect 169 -278 170 -274
rect 174 -278 175 -274
rect 177 -278 182 -274
rect 162 -282 166 -278
rect 158 -286 159 -282
rect 161 -286 166 -282
rect 146 -310 151 -306
rect 153 -310 154 -306
rect 146 -314 150 -310
rect 162 -290 166 -286
rect 178 -282 182 -278
rect 194 -266 198 -262
rect 236 -221 240 -219
rect 276 -217 280 -216
rect 373 -209 383 -208
rect 458 -209 462 -208
rect 401 -213 403 -209
rect 458 -212 462 -211
rect 393 -214 403 -213
rect 414 -216 498 -212
rect 502 -216 563 -212
rect 393 -217 403 -216
rect 426 -217 430 -216
rect 276 -221 280 -219
rect 236 -224 251 -221
rect 247 -225 251 -224
rect 268 -224 280 -221
rect 268 -225 272 -224
rect 426 -220 430 -219
rect 373 -222 383 -221
rect 247 -228 251 -227
rect 268 -228 272 -227
rect 247 -231 250 -228
rect 373 -225 383 -224
rect 442 -225 446 -224
rect 401 -229 403 -225
rect 442 -228 446 -227
rect 393 -230 403 -229
rect 414 -232 498 -228
rect 502 -232 563 -228
rect 393 -233 403 -232
rect 482 -233 486 -232
rect 538 -233 542 -232
rect 482 -236 486 -235
rect 538 -236 542 -235
rect 236 -249 240 -248
rect 236 -253 240 -251
rect 276 -249 280 -248
rect 276 -253 280 -251
rect 236 -256 251 -253
rect 247 -257 251 -256
rect 268 -256 280 -253
rect 268 -257 272 -256
rect 373 -254 383 -253
rect 194 -270 199 -266
rect 201 -270 202 -266
rect 247 -260 251 -259
rect 268 -260 272 -259
rect 247 -263 250 -260
rect 236 -265 240 -264
rect 194 -274 198 -270
rect 236 -269 240 -267
rect 276 -265 280 -264
rect 373 -257 383 -256
rect 426 -257 430 -256
rect 401 -261 403 -257
rect 426 -260 430 -259
rect 393 -262 403 -261
rect 414 -264 498 -260
rect 502 -264 563 -260
rect 393 -265 403 -264
rect 506 -265 510 -264
rect 538 -265 542 -264
rect 276 -269 280 -267
rect 236 -272 251 -269
rect 247 -273 251 -272
rect 194 -278 199 -274
rect 201 -278 202 -274
rect 268 -272 280 -269
rect 268 -273 272 -272
rect 506 -268 510 -267
rect 373 -270 383 -269
rect 538 -268 542 -267
rect 194 -282 198 -278
rect 178 -286 183 -282
rect 185 -286 186 -282
rect 190 -286 191 -282
rect 193 -286 198 -282
rect 178 -290 182 -286
rect 162 -294 167 -290
rect 169 -294 170 -290
rect 174 -294 175 -290
rect 177 -294 182 -290
rect 162 -306 166 -294
rect 162 -310 167 -306
rect 169 -310 170 -306
rect 162 -314 166 -310
rect 146 -318 151 -314
rect 153 -318 154 -314
rect 158 -318 159 -314
rect 161 -318 166 -314
rect 146 -322 150 -318
rect 130 -326 135 -322
rect 137 -326 138 -322
rect 142 -326 143 -322
rect 145 -326 150 -322
rect 130 -330 134 -326
rect 130 -334 135 -330
rect 137 -334 138 -330
rect 130 -338 134 -334
rect 146 -338 150 -326
rect 130 -342 135 -338
rect 137 -342 138 -338
rect 142 -342 143 -338
rect 145 -342 150 -338
rect 130 -346 134 -342
rect 130 -350 135 -346
rect 137 -350 138 -346
rect 130 -354 134 -350
rect 146 -354 150 -342
rect 130 -358 135 -354
rect 137 -358 138 -354
rect 142 -358 143 -354
rect 145 -358 150 -354
rect 130 -361 134 -358
rect 146 -361 150 -358
rect 162 -330 166 -318
rect 158 -334 159 -330
rect 161 -334 166 -330
rect 162 -338 166 -334
rect 162 -342 167 -338
rect 169 -342 170 -338
rect 162 -361 166 -342
rect 178 -298 182 -294
rect 194 -290 198 -286
rect 190 -294 191 -290
rect 193 -294 198 -290
rect 178 -302 183 -298
rect 185 -302 186 -298
rect 178 -306 182 -302
rect 178 -310 183 -306
rect 185 -310 186 -306
rect 178 -322 182 -310
rect 194 -298 198 -294
rect 247 -276 251 -275
rect 268 -276 272 -275
rect 247 -279 250 -276
rect 236 -281 240 -280
rect 236 -285 240 -283
rect 276 -281 280 -280
rect 373 -273 383 -272
rect 426 -273 430 -272
rect 401 -277 403 -273
rect 426 -276 430 -275
rect 393 -278 403 -277
rect 414 -280 498 -276
rect 502 -280 563 -276
rect 393 -281 403 -280
rect 426 -281 430 -280
rect 434 -281 438 -280
rect 276 -285 280 -283
rect 236 -288 251 -285
rect 247 -289 251 -288
rect 268 -288 280 -285
rect 268 -289 272 -288
rect 426 -284 430 -283
rect 373 -286 383 -285
rect 434 -284 438 -283
rect 194 -302 199 -298
rect 201 -302 202 -298
rect 247 -292 251 -291
rect 268 -292 272 -291
rect 247 -295 250 -292
rect 236 -297 240 -296
rect 194 -314 198 -302
rect 190 -318 191 -314
rect 193 -318 198 -314
rect 178 -326 183 -322
rect 185 -326 186 -322
rect 178 -346 182 -326
rect 174 -350 175 -346
rect 177 -350 182 -346
rect 178 -361 182 -350
rect 194 -330 198 -318
rect 236 -301 240 -299
rect 276 -297 280 -296
rect 373 -289 383 -288
rect 434 -289 438 -288
rect 401 -293 403 -289
rect 434 -292 438 -291
rect 393 -294 403 -293
rect 414 -296 498 -292
rect 502 -296 563 -292
rect 393 -297 403 -296
rect 458 -297 462 -296
rect 276 -301 280 -299
rect 236 -304 251 -301
rect 247 -305 251 -304
rect 268 -304 280 -301
rect 268 -305 272 -304
rect 458 -300 462 -299
rect 373 -302 383 -301
rect 247 -308 251 -307
rect 268 -308 272 -307
rect 247 -311 250 -308
rect 236 -313 240 -312
rect 236 -317 240 -315
rect 276 -313 280 -312
rect 373 -305 383 -304
rect 546 -305 550 -304
rect 401 -309 403 -305
rect 546 -308 550 -307
rect 393 -310 403 -309
rect 414 -312 498 -308
rect 502 -312 563 -308
rect 393 -313 403 -312
rect 538 -313 542 -312
rect 554 -313 558 -312
rect 276 -317 280 -315
rect 236 -320 251 -317
rect 247 -321 251 -320
rect 268 -320 280 -317
rect 268 -321 272 -320
rect 538 -316 542 -315
rect 373 -318 383 -317
rect 554 -316 558 -315
rect 194 -334 199 -330
rect 201 -334 202 -330
rect 247 -324 251 -323
rect 268 -324 272 -323
rect 247 -327 250 -324
rect 236 -329 240 -328
rect 194 -346 198 -334
rect 236 -333 240 -331
rect 276 -329 280 -328
rect 373 -321 383 -320
rect 442 -321 446 -320
rect 401 -325 403 -321
rect 442 -324 446 -323
rect 393 -326 403 -325
rect 414 -328 498 -324
rect 502 -328 563 -324
rect 393 -329 403 -328
rect 434 -329 438 -328
rect 276 -333 280 -331
rect 236 -336 251 -333
rect 247 -337 251 -336
rect 268 -336 280 -333
rect 268 -337 272 -336
rect 434 -332 438 -331
rect 373 -334 383 -333
rect 194 -350 199 -346
rect 201 -350 202 -346
rect 247 -340 251 -339
rect 268 -340 272 -339
rect 247 -343 250 -340
rect 276 -345 280 -344
rect 373 -337 383 -336
rect 442 -337 446 -336
rect 401 -341 403 -337
rect 442 -340 446 -339
rect 393 -342 403 -341
rect 414 -344 498 -340
rect 502 -344 563 -340
rect 393 -345 403 -344
rect 418 -345 422 -344
rect 276 -349 280 -347
rect 194 -354 198 -350
rect 194 -358 199 -354
rect 201 -358 202 -354
rect 268 -352 280 -349
rect 268 -353 272 -352
rect 418 -348 422 -347
rect 373 -350 383 -349
rect 268 -356 272 -355
rect 194 -361 198 -358
rect 373 -353 383 -352
rect 418 -353 422 -352
rect 442 -353 446 -352
rect 418 -356 422 -355
rect 442 -356 446 -355
rect 414 -360 498 -356
rect 502 -360 563 -356
rect 34 -380 37 -378
rect 36 -391 37 -380
rect 39 -391 40 -378
rect 50 -380 53 -378
rect 28 -415 29 -401
rect 31 -415 32 -401
rect 52 -391 53 -380
rect 55 -391 56 -378
rect 66 -380 69 -378
rect 44 -415 45 -401
rect 47 -415 48 -401
rect 68 -391 69 -380
rect 71 -391 72 -378
rect 82 -380 85 -378
rect 60 -415 61 -401
rect 63 -415 64 -401
rect 84 -391 85 -380
rect 87 -391 88 -378
rect 98 -380 101 -378
rect 76 -415 77 -401
rect 79 -415 80 -401
rect 100 -391 101 -380
rect 103 -391 104 -378
rect 114 -380 117 -378
rect 92 -415 93 -401
rect 95 -415 96 -401
rect 116 -391 117 -380
rect 119 -391 120 -378
rect 130 -380 133 -378
rect 108 -415 109 -401
rect 111 -415 112 -401
rect 132 -391 133 -380
rect 135 -391 136 -378
rect 146 -380 149 -378
rect 124 -415 125 -401
rect 127 -415 128 -401
rect 148 -391 149 -380
rect 151 -391 152 -378
rect 162 -380 165 -378
rect 140 -415 141 -401
rect 143 -415 144 -401
rect 164 -391 165 -380
rect 167 -391 168 -378
rect 178 -380 181 -378
rect 156 -415 157 -401
rect 159 -415 160 -401
rect 180 -391 181 -380
rect 183 -391 184 -378
rect 194 -380 197 -378
rect 172 -415 173 -401
rect 175 -415 176 -401
rect 196 -391 197 -380
rect 199 -391 200 -378
rect 427 -388 431 -376
rect 433 -383 434 -376
rect 433 -388 437 -383
rect 427 -391 430 -388
rect 188 -415 189 -401
rect 191 -415 192 -401
rect 419 -393 423 -391
rect 422 -403 423 -393
rect 425 -403 430 -391
rect 443 -388 447 -376
rect 449 -383 450 -376
rect 449 -388 453 -383
rect 443 -391 446 -388
rect 435 -393 439 -391
rect 438 -403 439 -393
rect 441 -403 446 -391
rect 459 -388 463 -376
rect 465 -383 466 -376
rect 465 -388 469 -383
rect 459 -391 462 -388
rect 451 -393 455 -391
rect 454 -403 455 -393
rect 457 -403 462 -391
rect 422 -553 423 -543
rect 38 -561 42 -560
rect 54 -561 58 -560
rect 70 -561 74 -560
rect 86 -561 90 -560
rect 102 -561 106 -560
rect 118 -561 122 -560
rect 134 -561 138 -560
rect 150 -561 154 -560
rect 166 -561 170 -560
rect 182 -561 186 -560
rect 419 -555 423 -553
rect 425 -555 430 -543
rect 427 -558 430 -555
rect 475 -388 479 -376
rect 481 -383 482 -376
rect 481 -388 485 -383
rect 475 -391 478 -388
rect 467 -393 471 -391
rect 470 -403 471 -393
rect 473 -403 478 -391
rect 438 -553 439 -543
rect 435 -555 439 -553
rect 441 -555 446 -543
rect 198 -561 202 -560
rect 38 -566 42 -563
rect 54 -566 58 -563
rect 70 -566 74 -563
rect 86 -566 90 -563
rect 102 -566 106 -563
rect 118 -566 122 -563
rect 134 -566 138 -563
rect 150 -566 154 -563
rect 166 -566 170 -563
rect 182 -566 186 -563
rect 198 -566 202 -563
rect 38 -569 42 -568
rect 54 -569 58 -568
rect 70 -569 74 -568
rect 86 -569 90 -568
rect 102 -569 106 -568
rect 118 -569 122 -568
rect 134 -569 138 -568
rect 150 -569 154 -568
rect 166 -569 170 -568
rect 182 -569 186 -568
rect 198 -569 202 -568
rect 427 -570 431 -558
rect 433 -563 437 -558
rect 443 -558 446 -555
rect 491 -388 495 -376
rect 497 -383 498 -376
rect 497 -388 501 -383
rect 491 -391 494 -388
rect 483 -393 487 -391
rect 486 -403 487 -393
rect 489 -403 494 -391
rect 454 -553 455 -543
rect 451 -555 455 -553
rect 457 -555 462 -543
rect 433 -570 434 -563
rect 443 -570 447 -558
rect 449 -563 453 -558
rect 459 -558 462 -555
rect 515 -388 519 -376
rect 521 -383 522 -376
rect 521 -388 525 -383
rect 515 -391 518 -388
rect 507 -393 511 -391
rect 510 -403 511 -393
rect 513 -403 518 -391
rect 470 -553 471 -543
rect 467 -555 471 -553
rect 473 -555 478 -543
rect 449 -570 450 -563
rect 459 -570 463 -558
rect 465 -563 469 -558
rect 475 -558 478 -555
rect 531 -388 535 -376
rect 537 -383 538 -376
rect 537 -388 541 -383
rect 531 -391 534 -388
rect 523 -393 527 -391
rect 526 -403 527 -393
rect 529 -403 534 -391
rect 486 -553 487 -543
rect 483 -555 487 -553
rect 489 -555 494 -543
rect 465 -570 466 -563
rect 475 -570 479 -558
rect 481 -563 485 -558
rect 491 -558 494 -555
rect 547 -388 551 -376
rect 553 -383 554 -376
rect 553 -388 557 -383
rect 547 -391 550 -388
rect 539 -393 543 -391
rect 542 -403 543 -393
rect 545 -403 550 -391
rect 510 -553 511 -543
rect 507 -555 511 -553
rect 513 -555 518 -543
rect 481 -570 482 -563
rect 491 -570 495 -558
rect 497 -563 501 -558
rect 515 -558 518 -555
rect 526 -553 527 -543
rect 523 -555 527 -553
rect 529 -555 534 -543
rect 497 -570 498 -563
rect 515 -570 519 -558
rect 521 -563 525 -558
rect 531 -558 534 -555
rect 542 -553 543 -543
rect 539 -555 543 -553
rect 545 -555 550 -543
rect 521 -570 522 -563
rect 531 -570 535 -558
rect 537 -563 541 -558
rect 547 -558 550 -555
rect 558 -553 559 -543
rect 555 -555 559 -553
rect 561 -555 566 -543
rect 537 -570 538 -563
rect 547 -570 551 -558
rect 553 -563 557 -558
rect 563 -558 566 -555
rect 553 -570 554 -563
rect 563 -570 567 -558
rect 569 -563 573 -558
rect 569 -570 570 -563
<< pdiffusion >>
rect 418 21 422 22
rect 426 21 430 22
rect 434 21 438 22
rect 442 21 446 22
rect 450 21 454 22
rect 458 21 462 22
rect 466 21 470 22
rect 474 21 478 22
rect 482 21 486 22
rect 490 21 494 22
rect 506 21 510 22
rect 514 21 518 22
rect 522 21 526 22
rect 530 21 534 22
rect 538 21 542 22
rect 546 21 550 22
rect 554 21 558 22
rect 418 18 422 19
rect 426 18 430 19
rect 434 18 438 19
rect 442 18 446 19
rect 450 18 454 19
rect 458 18 462 19
rect 466 18 470 19
rect 474 18 478 19
rect 482 18 486 19
rect 490 18 494 19
rect 506 18 510 19
rect 514 18 518 19
rect 522 18 526 19
rect 530 18 534 19
rect 538 18 542 19
rect 546 18 550 19
rect 554 18 558 19
rect 8 -6 9 -2
rect 11 -6 12 -2
rect 8 -14 9 -10
rect 11 -14 12 -10
rect 8 -22 9 -18
rect 11 -22 12 -18
rect 8 -30 9 -26
rect 11 -30 12 -26
rect 8 -38 9 -34
rect 11 -38 12 -34
rect 8 -46 9 -42
rect 11 -46 12 -42
rect 8 -54 9 -50
rect 11 -54 12 -50
rect 8 -62 9 -58
rect 11 -62 12 -58
rect 8 -70 9 -66
rect 11 -70 12 -66
rect 8 -78 9 -74
rect 11 -78 12 -74
rect 8 -86 9 -82
rect 11 -86 12 -82
rect 8 -94 9 -90
rect 11 -94 12 -90
rect 8 -102 9 -98
rect 11 -102 12 -98
rect 8 -110 9 -106
rect 11 -110 12 -106
rect 8 -134 9 -130
rect 11 -134 12 -130
rect 8 -142 9 -138
rect 11 -142 12 -138
rect 8 -150 9 -146
rect 11 -150 12 -146
rect 8 -158 9 -154
rect 11 -158 12 -154
rect 8 -166 9 -162
rect 11 -166 12 -162
rect 8 -174 9 -170
rect 11 -174 12 -170
rect 8 -182 9 -178
rect 11 -182 12 -178
rect 8 -190 9 -186
rect 11 -190 12 -186
rect 8 -198 9 -194
rect 11 -198 12 -194
rect 8 -206 9 -202
rect 11 -206 12 -202
rect 8 -214 9 -210
rect 11 -214 12 -210
rect 8 -222 9 -218
rect 11 -222 12 -218
rect 8 -230 9 -226
rect 11 -230 12 -226
rect 8 -238 9 -234
rect 11 -238 12 -234
rect 8 -262 9 -258
rect 11 -262 12 -258
rect 8 -270 9 -266
rect 11 -270 12 -266
rect 8 -278 9 -274
rect 11 -278 12 -274
rect 8 -286 9 -282
rect 11 -286 12 -282
rect 8 -294 9 -290
rect 11 -294 12 -290
rect 8 -302 9 -298
rect 11 -302 12 -298
rect 8 -310 9 -306
rect 11 -310 12 -306
rect 8 -318 9 -314
rect 11 -318 12 -314
rect 8 -326 9 -322
rect 11 -326 12 -322
rect 8 -334 9 -330
rect 11 -334 12 -330
rect 8 -342 9 -338
rect 11 -342 12 -338
rect 8 -350 9 -346
rect 11 -350 12 -346
rect 8 -358 9 -354
rect 11 -358 12 -354
rect 222 7 226 8
rect 222 4 226 5
rect 290 7 294 8
rect 222 -1 226 0
rect 290 4 294 5
rect 290 -1 294 0
rect 343 3 348 7
rect 343 2 363 3
rect 343 -1 363 0
rect 222 -4 226 -3
rect 290 -4 294 -3
rect 222 -9 226 -8
rect 222 -12 226 -11
rect 313 -5 315 -1
rect 290 -9 294 -8
rect 313 -6 333 -5
rect 313 -9 333 -8
rect 222 -17 226 -16
rect 290 -12 294 -11
rect 290 -17 294 -16
rect 313 -13 315 -9
rect 343 -13 348 -9
rect 343 -14 363 -13
rect 343 -17 363 -16
rect 222 -20 226 -19
rect 290 -20 294 -19
rect 222 -25 226 -24
rect 222 -28 226 -27
rect 313 -21 315 -17
rect 290 -25 294 -24
rect 313 -22 333 -21
rect 313 -25 333 -24
rect 222 -33 226 -32
rect 290 -28 294 -27
rect 290 -33 294 -32
rect 313 -29 315 -25
rect 343 -29 348 -25
rect 343 -30 363 -29
rect 343 -33 363 -32
rect 222 -36 226 -35
rect 290 -36 294 -35
rect 222 -41 226 -40
rect 222 -44 226 -43
rect 313 -37 315 -33
rect 290 -41 294 -40
rect 313 -38 333 -37
rect 313 -41 333 -40
rect 222 -49 226 -48
rect 290 -44 294 -43
rect 290 -49 294 -48
rect 313 -45 315 -41
rect 343 -45 348 -41
rect 343 -46 363 -45
rect 343 -49 363 -48
rect 222 -52 226 -51
rect 290 -52 294 -51
rect 222 -57 226 -56
rect 222 -60 226 -59
rect 313 -53 315 -49
rect 290 -57 294 -56
rect 313 -54 333 -53
rect 313 -57 333 -56
rect 222 -65 226 -64
rect 290 -60 294 -59
rect 290 -65 294 -64
rect 313 -61 315 -57
rect 343 -61 348 -57
rect 343 -62 363 -61
rect 343 -65 363 -64
rect 222 -68 226 -67
rect 290 -68 294 -67
rect 222 -73 226 -72
rect 222 -76 226 -75
rect 313 -69 315 -65
rect 290 -73 294 -72
rect 313 -70 333 -69
rect 313 -73 333 -72
rect 222 -81 226 -80
rect 290 -76 294 -75
rect 290 -81 294 -80
rect 313 -77 315 -73
rect 343 -77 348 -73
rect 343 -78 363 -77
rect 343 -81 363 -80
rect 222 -84 226 -83
rect 290 -84 294 -83
rect 222 -89 226 -88
rect 222 -92 226 -91
rect 313 -85 315 -81
rect 290 -89 294 -88
rect 313 -86 333 -85
rect 313 -89 333 -88
rect 222 -97 226 -96
rect 290 -92 294 -91
rect 290 -97 294 -96
rect 313 -93 315 -89
rect 343 -93 348 -89
rect 343 -94 363 -93
rect 343 -97 363 -96
rect 222 -100 226 -99
rect 290 -100 294 -99
rect 313 -101 315 -97
rect 313 -102 333 -101
rect 313 -105 333 -104
rect 313 -109 315 -105
rect 222 -121 226 -120
rect 222 -124 226 -123
rect 290 -121 294 -120
rect 222 -129 226 -128
rect 290 -124 294 -123
rect 290 -129 294 -128
rect 343 -125 348 -121
rect 343 -126 363 -125
rect 343 -129 363 -128
rect 222 -132 226 -131
rect 290 -132 294 -131
rect 222 -137 226 -136
rect 222 -140 226 -139
rect 313 -133 315 -129
rect 290 -137 294 -136
rect 313 -134 333 -133
rect 313 -137 333 -136
rect 222 -145 226 -144
rect 290 -140 294 -139
rect 290 -145 294 -144
rect 313 -141 315 -137
rect 343 -141 348 -137
rect 343 -142 363 -141
rect 343 -145 363 -144
rect 222 -148 226 -147
rect 290 -148 294 -147
rect 222 -153 226 -152
rect 222 -156 226 -155
rect 313 -149 315 -145
rect 290 -153 294 -152
rect 313 -150 333 -149
rect 313 -153 333 -152
rect 222 -161 226 -160
rect 290 -156 294 -155
rect 290 -161 294 -160
rect 313 -157 315 -153
rect 343 -157 348 -153
rect 343 -158 363 -157
rect 343 -161 363 -160
rect 222 -164 226 -163
rect 290 -164 294 -163
rect 222 -169 226 -168
rect 222 -172 226 -171
rect 313 -165 315 -161
rect 290 -169 294 -168
rect 313 -166 333 -165
rect 313 -169 333 -168
rect 222 -177 226 -176
rect 290 -172 294 -171
rect 290 -177 294 -176
rect 313 -173 315 -169
rect 343 -173 348 -169
rect 343 -174 363 -173
rect 343 -177 363 -176
rect 222 -180 226 -179
rect 290 -180 294 -179
rect 222 -185 226 -184
rect 222 -188 226 -187
rect 313 -181 315 -177
rect 290 -185 294 -184
rect 313 -182 333 -181
rect 313 -185 333 -184
rect 222 -193 226 -192
rect 290 -188 294 -187
rect 290 -193 294 -192
rect 313 -189 315 -185
rect 343 -189 348 -185
rect 343 -190 363 -189
rect 343 -193 363 -192
rect 222 -196 226 -195
rect 290 -196 294 -195
rect 222 -201 226 -200
rect 222 -204 226 -203
rect 313 -197 315 -193
rect 290 -201 294 -200
rect 313 -198 333 -197
rect 313 -201 333 -200
rect 222 -209 226 -208
rect 290 -204 294 -203
rect 290 -209 294 -208
rect 313 -205 315 -201
rect 343 -205 348 -201
rect 343 -206 363 -205
rect 343 -209 363 -208
rect 222 -212 226 -211
rect 290 -212 294 -211
rect 222 -217 226 -216
rect 222 -220 226 -219
rect 313 -213 315 -209
rect 290 -217 294 -216
rect 313 -214 333 -213
rect 313 -217 333 -216
rect 222 -225 226 -224
rect 290 -220 294 -219
rect 290 -225 294 -224
rect 313 -221 315 -217
rect 343 -221 348 -217
rect 343 -222 363 -221
rect 343 -225 363 -224
rect 222 -228 226 -227
rect 290 -228 294 -227
rect 313 -229 315 -225
rect 313 -230 333 -229
rect 313 -233 333 -232
rect 313 -237 315 -233
rect 222 -249 226 -248
rect 222 -252 226 -251
rect 290 -249 294 -248
rect 222 -257 226 -256
rect 290 -252 294 -251
rect 290 -257 294 -256
rect 343 -253 348 -249
rect 343 -254 363 -253
rect 343 -257 363 -256
rect 222 -260 226 -259
rect 290 -260 294 -259
rect 222 -265 226 -264
rect 222 -268 226 -267
rect 313 -261 315 -257
rect 290 -265 294 -264
rect 313 -262 333 -261
rect 313 -265 333 -264
rect 222 -273 226 -272
rect 290 -268 294 -267
rect 290 -273 294 -272
rect 313 -269 315 -265
rect 343 -269 348 -265
rect 343 -270 363 -269
rect 343 -273 363 -272
rect 222 -276 226 -275
rect 290 -276 294 -275
rect 222 -281 226 -280
rect 222 -284 226 -283
rect 313 -277 315 -273
rect 290 -281 294 -280
rect 313 -278 333 -277
rect 313 -281 333 -280
rect 222 -289 226 -288
rect 290 -284 294 -283
rect 290 -289 294 -288
rect 313 -285 315 -281
rect 343 -285 348 -281
rect 343 -286 363 -285
rect 343 -289 363 -288
rect 222 -292 226 -291
rect 290 -292 294 -291
rect 222 -297 226 -296
rect 222 -300 226 -299
rect 313 -293 315 -289
rect 290 -297 294 -296
rect 313 -294 333 -293
rect 313 -297 333 -296
rect 222 -305 226 -304
rect 290 -300 294 -299
rect 290 -305 294 -304
rect 313 -301 315 -297
rect 343 -301 348 -297
rect 343 -302 363 -301
rect 343 -305 363 -304
rect 222 -308 226 -307
rect 290 -308 294 -307
rect 222 -313 226 -312
rect 222 -316 226 -315
rect 313 -309 315 -305
rect 290 -313 294 -312
rect 313 -310 333 -309
rect 313 -313 333 -312
rect 222 -321 226 -320
rect 290 -316 294 -315
rect 290 -321 294 -320
rect 313 -317 315 -313
rect 343 -317 348 -313
rect 343 -318 363 -317
rect 343 -321 363 -320
rect 222 -324 226 -323
rect 290 -324 294 -323
rect 222 -329 226 -328
rect 222 -332 226 -331
rect 313 -325 315 -321
rect 290 -329 294 -328
rect 313 -326 333 -325
rect 313 -329 333 -328
rect 222 -337 226 -336
rect 290 -332 294 -331
rect 290 -337 294 -336
rect 313 -333 315 -329
rect 343 -333 348 -329
rect 343 -334 363 -333
rect 343 -337 363 -336
rect 222 -340 226 -339
rect 290 -340 294 -339
rect 313 -341 315 -337
rect 290 -345 294 -344
rect 313 -342 333 -341
rect 313 -345 333 -344
rect 290 -348 294 -347
rect 290 -353 294 -352
rect 313 -349 315 -345
rect 343 -349 348 -345
rect 343 -350 363 -349
rect 343 -353 363 -352
rect 290 -356 294 -355
rect 28 -444 29 -425
rect 26 -451 29 -444
rect 31 -451 32 -425
rect 44 -444 45 -425
rect 42 -451 45 -444
rect 47 -451 48 -425
rect 36 -485 37 -461
rect 32 -487 37 -485
rect 39 -478 40 -461
rect 39 -487 42 -478
rect 60 -444 61 -425
rect 58 -451 61 -444
rect 63 -451 64 -425
rect 52 -485 53 -461
rect 48 -487 53 -485
rect 55 -478 56 -461
rect 55 -487 58 -478
rect 76 -444 77 -425
rect 74 -451 77 -444
rect 79 -451 80 -425
rect 68 -485 69 -461
rect 64 -487 69 -485
rect 71 -478 72 -461
rect 71 -487 74 -478
rect 92 -444 93 -425
rect 90 -451 93 -444
rect 95 -451 96 -425
rect 84 -485 85 -461
rect 80 -487 85 -485
rect 87 -478 88 -461
rect 87 -487 90 -478
rect 108 -444 109 -425
rect 106 -451 109 -444
rect 111 -451 112 -425
rect 100 -485 101 -461
rect 96 -487 101 -485
rect 103 -478 104 -461
rect 103 -487 106 -478
rect 124 -444 125 -425
rect 122 -451 125 -444
rect 127 -451 128 -425
rect 116 -485 117 -461
rect 112 -487 117 -485
rect 119 -478 120 -461
rect 119 -487 122 -478
rect 140 -444 141 -425
rect 138 -451 141 -444
rect 143 -451 144 -425
rect 132 -485 133 -461
rect 128 -487 133 -485
rect 135 -478 136 -461
rect 135 -487 138 -478
rect 156 -444 157 -425
rect 154 -451 157 -444
rect 159 -451 160 -425
rect 148 -485 149 -461
rect 144 -487 149 -485
rect 151 -478 152 -461
rect 151 -487 154 -478
rect 172 -444 173 -425
rect 170 -451 173 -444
rect 175 -451 176 -425
rect 164 -485 165 -461
rect 160 -487 165 -485
rect 167 -478 168 -461
rect 167 -487 170 -478
rect 188 -444 189 -425
rect 186 -451 189 -444
rect 191 -451 192 -425
rect 180 -485 181 -461
rect 176 -487 181 -485
rect 183 -478 184 -461
rect 183 -487 186 -478
rect 422 -435 423 -413
rect 419 -437 423 -435
rect 425 -437 430 -413
rect 427 -440 430 -437
rect 438 -435 439 -413
rect 435 -437 439 -435
rect 441 -437 446 -413
rect 196 -485 197 -461
rect 192 -487 197 -485
rect 199 -478 200 -461
rect 199 -487 202 -478
rect 38 -503 42 -502
rect 54 -503 58 -502
rect 70 -503 74 -502
rect 86 -503 90 -502
rect 102 -503 106 -502
rect 118 -503 122 -502
rect 134 -503 138 -502
rect 150 -503 154 -502
rect 166 -503 170 -502
rect 182 -503 186 -502
rect 198 -503 202 -502
rect 38 -508 42 -505
rect 54 -508 58 -505
rect 70 -508 74 -505
rect 86 -508 90 -505
rect 102 -508 106 -505
rect 118 -508 122 -505
rect 134 -508 138 -505
rect 150 -508 154 -505
rect 166 -508 170 -505
rect 182 -508 186 -505
rect 198 -508 202 -505
rect 427 -464 431 -440
rect 433 -445 437 -440
rect 443 -440 446 -437
rect 454 -435 455 -413
rect 451 -437 455 -435
rect 457 -437 462 -413
rect 433 -464 434 -445
rect 427 -505 431 -481
rect 433 -505 434 -481
rect 427 -509 430 -505
rect 38 -511 42 -510
rect 54 -511 58 -510
rect 70 -511 74 -510
rect 86 -511 90 -510
rect 102 -511 106 -510
rect 118 -511 122 -510
rect 134 -511 138 -510
rect 150 -511 154 -510
rect 166 -511 170 -510
rect 182 -511 186 -510
rect 198 -511 202 -510
rect 38 -534 42 -533
rect 54 -534 58 -533
rect 70 -534 74 -533
rect 86 -534 90 -533
rect 102 -534 106 -533
rect 118 -534 122 -533
rect 134 -534 138 -533
rect 150 -534 154 -533
rect 166 -534 170 -533
rect 182 -534 186 -533
rect 422 -533 423 -509
rect 425 -533 430 -509
rect 198 -534 202 -533
rect 38 -539 42 -536
rect 54 -539 58 -536
rect 70 -539 74 -536
rect 86 -539 90 -536
rect 102 -539 106 -536
rect 118 -539 122 -536
rect 134 -539 138 -536
rect 150 -539 154 -536
rect 166 -539 170 -536
rect 182 -539 186 -536
rect 198 -539 202 -536
rect 38 -542 42 -541
rect 54 -542 58 -541
rect 70 -542 74 -541
rect 86 -542 90 -541
rect 102 -542 106 -541
rect 118 -542 122 -541
rect 134 -542 138 -541
rect 150 -542 154 -541
rect 166 -542 170 -541
rect 182 -542 186 -541
rect 198 -542 202 -541
rect 443 -464 447 -440
rect 449 -445 453 -440
rect 459 -440 462 -437
rect 470 -435 471 -413
rect 467 -437 471 -435
rect 473 -437 478 -413
rect 449 -464 450 -445
rect 443 -505 447 -481
rect 449 -505 450 -481
rect 443 -509 446 -505
rect 438 -533 439 -509
rect 441 -533 446 -509
rect 459 -464 463 -440
rect 465 -445 469 -440
rect 475 -440 478 -437
rect 486 -435 487 -413
rect 483 -437 487 -435
rect 489 -437 494 -413
rect 465 -464 466 -445
rect 459 -505 463 -481
rect 465 -505 466 -481
rect 459 -509 462 -505
rect 454 -533 455 -509
rect 457 -533 462 -509
rect 475 -464 479 -440
rect 481 -445 485 -440
rect 491 -440 494 -437
rect 510 -435 511 -413
rect 507 -437 511 -435
rect 513 -437 518 -413
rect 481 -464 482 -445
rect 475 -505 479 -481
rect 481 -505 482 -481
rect 475 -509 478 -505
rect 470 -533 471 -509
rect 473 -533 478 -509
rect 491 -464 495 -440
rect 497 -445 501 -440
rect 515 -440 518 -437
rect 526 -435 527 -413
rect 523 -437 527 -435
rect 529 -437 534 -413
rect 497 -464 498 -445
rect 491 -505 495 -481
rect 497 -505 498 -481
rect 491 -509 494 -505
rect 486 -533 487 -509
rect 489 -533 494 -509
rect 515 -464 519 -440
rect 521 -445 525 -440
rect 531 -440 534 -437
rect 542 -435 543 -413
rect 539 -437 543 -435
rect 545 -437 550 -413
rect 521 -464 522 -445
rect 515 -505 519 -481
rect 521 -505 522 -481
rect 515 -509 518 -505
rect 510 -533 511 -509
rect 513 -533 518 -509
rect 531 -464 535 -440
rect 537 -445 541 -440
rect 547 -440 550 -437
rect 537 -464 538 -445
rect 531 -505 535 -481
rect 537 -505 538 -481
rect 531 -509 534 -505
rect 526 -533 527 -509
rect 529 -533 534 -509
rect 547 -464 551 -440
rect 553 -445 557 -440
rect 553 -464 554 -445
rect 547 -505 551 -481
rect 553 -505 554 -481
rect 547 -509 550 -505
rect 542 -533 543 -509
rect 545 -533 550 -509
rect 563 -505 567 -481
rect 569 -505 570 -481
rect 563 -509 566 -505
rect 558 -533 559 -509
rect 561 -533 566 -509
<< metal1 >>
rect 15 26 26 30
rect 206 26 390 30
rect 15 24 390 26
rect 15 16 19 24
rect 254 12 258 24
rect 230 8 236 11
rect 244 8 247 12
rect 7 7 11 8
rect 27 2 34 5
rect 38 2 50 5
rect 54 2 66 5
rect 70 2 82 5
rect 86 2 98 5
rect 102 2 114 5
rect 118 2 130 5
rect 134 2 146 5
rect 150 2 162 5
rect 166 2 178 5
rect 182 2 194 5
rect 198 2 206 5
rect 16 -6 42 -3
rect 46 -6 106 -3
rect 110 -6 122 -3
rect 126 -6 154 -3
rect 158 -6 170 -3
rect 174 -6 186 -3
rect 190 -6 202 -3
rect 206 -6 207 -2
rect 215 -4 219 8
rect 230 4 233 8
rect 226 1 229 4
rect 230 -8 236 -5
rect 244 -8 247 4
rect 254 -4 258 8
rect 261 -4 265 -3
rect 268 -4 272 24
rect 297 13 379 17
rect 297 12 301 13
rect 280 8 286 11
rect 283 4 286 8
rect 287 1 290 4
rect 297 -4 301 8
rect 341 -1 345 13
rect 386 10 390 24
rect 413 22 416 26
rect 560 22 562 26
rect 405 15 409 18
rect 565 18 569 19
rect 363 4 373 7
rect 366 -1 369 4
rect 386 6 409 10
rect 386 -1 390 6
rect 418 4 421 14
rect 280 -8 286 -5
rect 408 -5 409 -1
rect 16 -14 42 -11
rect 46 -14 58 -11
rect 62 -14 138 -11
rect 142 -14 154 -11
rect 158 -14 170 -11
rect 174 -14 186 -11
rect 190 -14 202 -11
rect 206 -14 208 -10
rect 16 -22 42 -19
rect 46 -22 74 -19
rect 78 -22 138 -19
rect 142 -22 170 -19
rect 174 -22 202 -19
rect 206 -22 207 -18
rect 215 -20 219 -8
rect 230 -12 233 -8
rect 226 -15 229 -12
rect 230 -24 236 -21
rect 244 -24 247 -12
rect 254 -20 258 -8
rect 261 -20 265 -19
rect 268 -20 272 -8
rect 283 -12 286 -8
rect 287 -15 290 -12
rect 297 -20 301 -8
rect 333 -13 334 -9
rect 341 -17 345 -5
rect 363 -12 373 -9
rect 366 -17 369 -12
rect 386 -17 390 -5
rect 403 -13 404 -9
rect 408 -13 409 -9
rect 418 -12 421 0
rect 426 -12 429 14
rect 434 -12 437 14
rect 280 -24 286 -21
rect 408 -21 409 -17
rect 16 -30 42 -27
rect 46 -30 74 -27
rect 78 -30 154 -27
rect 158 -30 170 -27
rect 174 -30 186 -27
rect 206 -27 208 -26
rect 190 -30 208 -27
rect 16 -38 42 -35
rect 46 -38 58 -35
rect 62 -38 138 -35
rect 142 -38 170 -35
rect 174 -38 186 -35
rect 206 -35 207 -34
rect 190 -38 207 -35
rect 215 -36 219 -24
rect 230 -28 233 -24
rect 226 -31 229 -28
rect 230 -40 236 -37
rect 244 -40 247 -28
rect 254 -36 258 -24
rect 261 -36 265 -35
rect 268 -36 272 -24
rect 283 -28 286 -24
rect 287 -31 290 -28
rect 297 -36 301 -24
rect 333 -29 334 -25
rect 341 -33 345 -21
rect 363 -28 373 -25
rect 366 -33 369 -28
rect 386 -33 390 -21
rect 403 -29 404 -25
rect 408 -29 409 -25
rect 418 -28 421 -16
rect 280 -40 286 -37
rect 408 -37 409 -33
rect 16 -46 42 -43
rect 46 -46 122 -43
rect 126 -46 154 -43
rect 158 -46 170 -43
rect 174 -46 202 -43
rect 206 -46 208 -42
rect 16 -54 42 -51
rect 46 -54 90 -51
rect 94 -54 122 -51
rect 126 -54 154 -51
rect 158 -54 170 -51
rect 174 -54 202 -51
rect 206 -54 207 -50
rect 215 -52 219 -40
rect 230 -44 233 -40
rect 226 -47 229 -44
rect 230 -56 236 -53
rect 244 -56 247 -44
rect 254 -52 258 -40
rect 261 -52 265 -51
rect 268 -52 272 -40
rect 283 -44 286 -40
rect 287 -47 290 -44
rect 297 -52 301 -40
rect 333 -45 334 -41
rect 341 -49 345 -37
rect 363 -44 373 -41
rect 366 -49 369 -44
rect 386 -49 390 -37
rect 403 -45 404 -41
rect 408 -45 409 -41
rect 280 -56 286 -53
rect 408 -53 409 -49
rect 16 -62 42 -59
rect 46 -62 90 -59
rect 94 -62 122 -59
rect 126 -62 154 -59
rect 158 -62 186 -59
rect 206 -59 208 -58
rect 190 -62 208 -59
rect 16 -70 42 -67
rect 46 -70 138 -67
rect 142 -70 154 -67
rect 158 -70 170 -67
rect 174 -70 186 -67
rect 206 -67 207 -66
rect 190 -70 207 -67
rect 215 -68 219 -56
rect 230 -60 233 -56
rect 226 -63 229 -60
rect 230 -72 236 -69
rect 244 -72 247 -60
rect 254 -68 258 -56
rect 261 -68 265 -67
rect 268 -68 272 -56
rect 283 -60 286 -56
rect 287 -63 290 -60
rect 297 -68 301 -56
rect 333 -61 334 -57
rect 341 -65 345 -53
rect 363 -60 373 -57
rect 366 -65 369 -60
rect 386 -65 390 -53
rect 403 -61 404 -57
rect 408 -61 409 -57
rect 418 -60 421 -32
rect 426 -44 429 -16
rect 434 -28 437 -16
rect 280 -72 286 -69
rect 408 -69 409 -65
rect 16 -78 42 -75
rect 46 -78 90 -75
rect 94 -78 122 -75
rect 126 -78 154 -75
rect 158 -78 170 -75
rect 206 -75 208 -74
rect 174 -78 208 -75
rect 16 -86 42 -83
rect 46 -86 122 -83
rect 126 -86 154 -83
rect 158 -86 186 -83
rect 190 -86 202 -83
rect 206 -86 207 -82
rect 215 -84 219 -72
rect 230 -76 233 -72
rect 226 -79 229 -76
rect 230 -88 236 -85
rect 244 -88 247 -76
rect 254 -84 258 -72
rect 261 -84 265 -83
rect 268 -84 272 -72
rect 283 -76 286 -72
rect 287 -79 290 -76
rect 297 -84 301 -72
rect 333 -77 334 -73
rect 341 -81 345 -69
rect 363 -76 373 -73
rect 366 -81 369 -76
rect 386 -81 390 -69
rect 403 -77 404 -73
rect 408 -77 409 -73
rect 418 -76 421 -64
rect 426 -76 429 -48
rect 434 -60 437 -32
rect 434 -76 437 -64
rect 280 -88 286 -85
rect 408 -85 409 -81
rect 16 -94 122 -91
rect 126 -94 154 -91
rect 158 -94 186 -91
rect 206 -91 208 -90
rect 190 -94 208 -91
rect 16 -102 138 -99
rect 142 -102 154 -99
rect 158 -102 186 -99
rect 206 -99 207 -98
rect 190 -102 207 -99
rect 215 -100 219 -88
rect 230 -92 233 -88
rect 226 -95 229 -92
rect 16 -110 138 -107
rect 142 -110 154 -107
rect 158 -110 170 -107
rect 174 -110 186 -107
rect 206 -107 208 -106
rect 190 -110 208 -107
rect 27 -118 34 -115
rect 38 -118 50 -115
rect 54 -118 66 -115
rect 70 -118 82 -115
rect 86 -118 98 -115
rect 102 -118 114 -115
rect 118 -118 130 -115
rect 134 -118 146 -115
rect 150 -118 162 -115
rect 166 -118 178 -115
rect 182 -118 194 -115
rect 198 -118 206 -115
rect 215 -116 219 -104
rect 230 -120 236 -117
rect 244 -120 247 -92
rect 254 -100 258 -88
rect 261 -100 265 -99
rect 268 -100 272 -88
rect 283 -92 286 -88
rect 287 -95 290 -92
rect 297 -100 301 -88
rect 333 -93 334 -89
rect 341 -97 345 -85
rect 363 -92 373 -89
rect 366 -97 369 -92
rect 386 -97 390 -85
rect 403 -93 404 -89
rect 408 -93 409 -89
rect 408 -101 409 -97
rect 19 -126 26 -122
rect 30 -126 42 -122
rect 46 -126 58 -122
rect 62 -126 74 -122
rect 78 -126 90 -122
rect 94 -126 106 -122
rect 110 -126 122 -122
rect 126 -126 138 -122
rect 142 -126 154 -122
rect 158 -126 170 -122
rect 174 -126 186 -122
rect 190 -126 202 -122
rect 16 -134 138 -131
rect 142 -134 154 -131
rect 158 -134 170 -131
rect 174 -134 202 -131
rect 206 -134 207 -130
rect 215 -132 219 -120
rect 230 -124 233 -120
rect 226 -127 229 -124
rect 230 -136 236 -133
rect 244 -136 247 -124
rect 254 -116 258 -104
rect 254 -132 258 -120
rect 261 -132 265 -131
rect 268 -132 272 -104
rect 297 -116 301 -104
rect 333 -109 334 -105
rect 280 -120 286 -117
rect 283 -124 286 -120
rect 287 -127 290 -124
rect 297 -132 301 -120
rect 341 -129 345 -101
rect 386 -116 390 -101
rect 403 -109 404 -105
rect 408 -109 409 -105
rect 363 -124 373 -121
rect 366 -129 369 -124
rect 386 -129 390 -120
rect 280 -136 286 -133
rect 408 -133 409 -129
rect 16 -142 122 -139
rect 126 -142 154 -139
rect 158 -142 170 -139
rect 174 -142 186 -139
rect 206 -139 208 -138
rect 190 -142 208 -139
rect 16 -150 122 -147
rect 126 -150 154 -147
rect 158 -150 170 -147
rect 174 -150 186 -147
rect 206 -147 207 -146
rect 190 -150 207 -147
rect 215 -148 219 -136
rect 230 -140 233 -136
rect 226 -143 229 -140
rect 230 -152 236 -149
rect 244 -152 247 -140
rect 254 -148 258 -136
rect 261 -148 265 -147
rect 268 -148 272 -136
rect 283 -140 286 -136
rect 287 -143 290 -140
rect 297 -148 301 -136
rect 333 -141 334 -137
rect 341 -145 345 -133
rect 363 -140 373 -137
rect 366 -145 369 -140
rect 386 -145 390 -133
rect 403 -141 404 -137
rect 408 -141 409 -137
rect 280 -152 286 -149
rect 408 -149 409 -145
rect 16 -158 42 -155
rect 46 -158 58 -155
rect 62 -158 138 -155
rect 142 -158 154 -155
rect 158 -158 202 -155
rect 206 -158 208 -154
rect 16 -166 42 -163
rect 46 -166 138 -163
rect 142 -166 186 -163
rect 206 -163 207 -162
rect 190 -166 207 -163
rect 215 -164 219 -152
rect 230 -156 233 -152
rect 226 -159 229 -156
rect 230 -168 236 -165
rect 244 -168 247 -156
rect 254 -164 258 -152
rect 261 -164 265 -163
rect 268 -164 272 -152
rect 283 -156 286 -152
rect 287 -159 290 -156
rect 297 -164 301 -152
rect 333 -157 334 -153
rect 341 -161 345 -149
rect 363 -156 373 -153
rect 366 -161 369 -156
rect 386 -161 390 -149
rect 403 -157 404 -153
rect 408 -157 409 -153
rect 418 -156 421 -80
rect 426 -156 429 -80
rect 280 -168 286 -165
rect 408 -165 409 -161
rect 16 -174 42 -171
rect 46 -174 122 -171
rect 126 -174 154 -171
rect 158 -174 170 -171
rect 174 -174 186 -171
rect 206 -171 208 -170
rect 190 -174 208 -171
rect 16 -182 138 -179
rect 142 -182 154 -179
rect 158 -182 170 -179
rect 174 -182 202 -179
rect 206 -182 207 -178
rect 215 -180 219 -168
rect 230 -172 233 -168
rect 226 -175 229 -172
rect 230 -184 236 -181
rect 244 -184 247 -172
rect 254 -180 258 -168
rect 261 -180 265 -179
rect 268 -180 272 -168
rect 283 -172 286 -168
rect 287 -175 290 -172
rect 297 -180 301 -168
rect 333 -173 334 -169
rect 341 -177 345 -165
rect 363 -172 373 -169
rect 366 -177 369 -172
rect 386 -177 390 -165
rect 403 -173 404 -169
rect 408 -173 409 -169
rect 418 -172 421 -160
rect 280 -184 286 -181
rect 408 -181 409 -177
rect 16 -190 138 -187
rect 142 -190 170 -187
rect 174 -190 202 -187
rect 206 -190 208 -186
rect 16 -198 138 -195
rect 142 -198 170 -195
rect 174 -198 186 -195
rect 206 -195 207 -194
rect 190 -198 207 -195
rect 215 -196 219 -184
rect 230 -188 233 -184
rect 226 -191 229 -188
rect 230 -200 236 -197
rect 244 -200 247 -188
rect 254 -196 258 -184
rect 261 -196 265 -195
rect 268 -196 272 -184
rect 283 -188 286 -184
rect 287 -191 290 -188
rect 297 -196 301 -184
rect 333 -189 334 -185
rect 341 -193 345 -181
rect 363 -188 373 -185
rect 366 -193 369 -188
rect 386 -193 390 -181
rect 403 -189 404 -185
rect 408 -189 409 -185
rect 280 -200 286 -197
rect 408 -197 409 -193
rect 16 -206 42 -203
rect 46 -206 122 -203
rect 126 -206 154 -203
rect 158 -206 170 -203
rect 206 -203 208 -202
rect 174 -206 208 -203
rect 16 -214 138 -211
rect 142 -214 154 -211
rect 158 -214 170 -211
rect 174 -214 186 -211
rect 206 -211 207 -210
rect 190 -214 207 -211
rect 215 -212 219 -200
rect 230 -204 233 -200
rect 226 -207 229 -204
rect 230 -216 236 -213
rect 244 -216 247 -204
rect 254 -212 258 -200
rect 261 -212 265 -211
rect 268 -212 272 -200
rect 283 -204 286 -200
rect 287 -207 290 -204
rect 297 -212 301 -200
rect 333 -205 334 -201
rect 341 -209 345 -197
rect 363 -204 373 -201
rect 366 -209 369 -204
rect 386 -209 390 -197
rect 403 -205 404 -201
rect 408 -205 409 -201
rect 280 -216 286 -213
rect 408 -213 409 -209
rect 16 -222 42 -219
rect 46 -222 138 -219
rect 142 -222 170 -219
rect 174 -222 202 -219
rect 206 -222 208 -218
rect 16 -230 42 -227
rect 46 -230 138 -227
rect 142 -230 154 -227
rect 158 -230 170 -227
rect 206 -227 207 -226
rect 174 -230 207 -227
rect 215 -228 219 -216
rect 230 -220 233 -216
rect 226 -223 229 -220
rect 16 -238 138 -235
rect 142 -238 154 -235
rect 158 -238 170 -235
rect 174 -238 186 -235
rect 206 -235 208 -234
rect 190 -238 208 -235
rect 27 -246 34 -243
rect 38 -246 50 -243
rect 54 -246 66 -243
rect 70 -246 82 -243
rect 86 -246 98 -243
rect 102 -246 114 -243
rect 118 -246 130 -243
rect 134 -246 146 -243
rect 150 -246 162 -243
rect 166 -246 178 -243
rect 182 -246 194 -243
rect 198 -246 206 -243
rect 215 -244 219 -232
rect 230 -248 236 -245
rect 244 -248 247 -220
rect 254 -228 258 -216
rect 261 -228 265 -227
rect 268 -228 272 -216
rect 283 -220 286 -216
rect 287 -223 290 -220
rect 297 -228 301 -216
rect 333 -221 334 -217
rect 341 -225 345 -213
rect 363 -220 373 -217
rect 366 -225 369 -220
rect 386 -225 390 -213
rect 403 -221 404 -217
rect 408 -221 409 -217
rect 408 -229 409 -225
rect 19 -254 26 -250
rect 30 -254 42 -250
rect 46 -254 58 -250
rect 62 -254 74 -250
rect 78 -254 90 -250
rect 94 -254 106 -250
rect 110 -254 122 -250
rect 126 -254 138 -250
rect 142 -254 154 -250
rect 158 -254 170 -250
rect 174 -254 186 -250
rect 190 -254 202 -250
rect 16 -262 42 -259
rect 46 -262 154 -259
rect 158 -262 170 -259
rect 174 -262 186 -259
rect 206 -259 207 -258
rect 190 -262 207 -259
rect 215 -260 219 -248
rect 230 -252 233 -248
rect 226 -255 229 -252
rect 230 -264 236 -261
rect 244 -264 247 -252
rect 254 -244 258 -232
rect 254 -260 258 -248
rect 261 -260 265 -259
rect 268 -260 272 -232
rect 297 -244 301 -232
rect 333 -237 334 -233
rect 280 -248 286 -245
rect 283 -252 286 -248
rect 287 -255 290 -252
rect 297 -260 301 -248
rect 341 -257 345 -229
rect 386 -244 390 -229
rect 403 -237 404 -233
rect 408 -237 409 -233
rect 363 -252 373 -249
rect 366 -257 369 -252
rect 386 -257 390 -248
rect 280 -264 286 -261
rect 408 -261 409 -257
rect 16 -270 138 -267
rect 142 -270 154 -267
rect 158 -270 170 -267
rect 174 -270 202 -267
rect 206 -270 208 -266
rect 16 -278 42 -275
rect 46 -278 154 -275
rect 158 -278 170 -275
rect 174 -278 202 -275
rect 206 -278 207 -274
rect 215 -276 219 -264
rect 230 -268 233 -264
rect 226 -271 229 -268
rect 230 -280 236 -277
rect 244 -280 247 -268
rect 254 -276 258 -264
rect 261 -276 265 -275
rect 268 -276 272 -264
rect 283 -268 286 -264
rect 287 -271 290 -268
rect 297 -276 301 -264
rect 333 -269 334 -265
rect 341 -273 345 -261
rect 363 -268 373 -265
rect 366 -273 369 -268
rect 386 -273 390 -261
rect 403 -269 404 -265
rect 408 -269 409 -265
rect 280 -280 286 -277
rect 408 -277 409 -273
rect 16 -286 42 -283
rect 46 -286 138 -283
rect 142 -286 154 -283
rect 158 -286 186 -283
rect 206 -283 208 -282
rect 190 -286 208 -283
rect 16 -294 42 -291
rect 46 -294 138 -291
rect 142 -294 170 -291
rect 174 -294 186 -291
rect 206 -291 207 -290
rect 190 -294 207 -291
rect 215 -292 219 -280
rect 230 -284 233 -280
rect 226 -287 229 -284
rect 230 -296 236 -293
rect 244 -296 247 -284
rect 254 -292 258 -280
rect 261 -292 265 -291
rect 268 -292 272 -280
rect 283 -284 286 -280
rect 287 -287 290 -284
rect 297 -292 301 -280
rect 333 -285 334 -281
rect 341 -289 345 -277
rect 363 -284 373 -281
rect 366 -289 369 -284
rect 386 -289 390 -277
rect 403 -285 404 -281
rect 408 -285 409 -281
rect 280 -296 286 -293
rect 408 -293 409 -289
rect 16 -302 138 -299
rect 142 -302 186 -299
rect 190 -302 202 -299
rect 206 -302 208 -298
rect 16 -310 122 -307
rect 126 -310 154 -307
rect 158 -310 170 -307
rect 174 -310 186 -307
rect 206 -307 207 -306
rect 190 -310 207 -307
rect 215 -308 219 -296
rect 230 -300 233 -296
rect 226 -303 229 -300
rect 230 -312 236 -309
rect 244 -312 247 -300
rect 254 -308 258 -296
rect 261 -308 265 -307
rect 268 -308 272 -296
rect 283 -300 286 -296
rect 287 -303 290 -300
rect 297 -308 301 -296
rect 333 -301 334 -297
rect 341 -305 345 -293
rect 363 -300 373 -297
rect 366 -305 369 -300
rect 386 -305 390 -293
rect 403 -301 404 -297
rect 408 -301 409 -297
rect 280 -312 286 -309
rect 408 -309 409 -305
rect 16 -318 138 -315
rect 142 -318 154 -315
rect 158 -318 186 -315
rect 206 -315 208 -314
rect 190 -318 208 -315
rect 16 -326 42 -323
rect 46 -326 138 -323
rect 142 -326 186 -323
rect 206 -323 207 -322
rect 190 -326 207 -323
rect 215 -324 219 -312
rect 230 -316 233 -312
rect 226 -319 229 -316
rect 230 -328 236 -325
rect 244 -328 247 -316
rect 254 -324 258 -312
rect 261 -324 265 -323
rect 268 -324 272 -312
rect 283 -316 286 -312
rect 287 -319 290 -316
rect 297 -324 301 -312
rect 333 -317 334 -313
rect 341 -321 345 -309
rect 363 -316 373 -313
rect 366 -321 369 -316
rect 386 -321 390 -309
rect 403 -317 404 -313
rect 408 -317 409 -313
rect 280 -328 286 -325
rect 408 -325 409 -321
rect 16 -334 42 -331
rect 46 -334 138 -331
rect 142 -334 154 -331
rect 158 -334 202 -331
rect 206 -334 208 -330
rect 16 -342 42 -339
rect 46 -342 138 -339
rect 142 -342 170 -339
rect 206 -339 207 -338
rect 174 -342 207 -339
rect 215 -340 219 -328
rect 230 -332 233 -328
rect 226 -335 229 -332
rect 244 -344 247 -332
rect 254 -340 258 -328
rect 261 -340 265 -339
rect 268 -340 272 -328
rect 283 -332 286 -328
rect 287 -335 290 -332
rect 297 -340 301 -328
rect 333 -333 334 -329
rect 341 -337 345 -325
rect 363 -332 373 -329
rect 366 -337 369 -332
rect 386 -337 390 -325
rect 403 -333 404 -329
rect 408 -333 409 -329
rect 280 -344 286 -341
rect 408 -341 409 -337
rect 16 -350 42 -347
rect 46 -350 138 -347
rect 142 -350 170 -347
rect 174 -350 202 -347
rect 206 -350 208 -346
rect 16 -358 42 -355
rect 46 -358 138 -355
rect 142 -358 202 -355
rect 206 -358 207 -354
rect 215 -356 219 -344
rect 0 -481 4 -360
rect 27 -365 34 -362
rect 38 -365 50 -362
rect 54 -365 66 -362
rect 70 -365 82 -362
rect 86 -365 98 -362
rect 102 -365 114 -362
rect 118 -365 130 -362
rect 134 -365 146 -362
rect 150 -365 162 -362
rect 166 -365 178 -362
rect 182 -365 194 -362
rect 198 -365 212 -362
rect 215 -364 224 -360
rect 7 -368 11 -367
rect 0 -511 4 -485
rect 8 -503 11 -372
rect 32 -373 36 -372
rect 40 -373 44 -372
rect 48 -373 52 -372
rect 56 -373 60 -372
rect 64 -373 68 -372
rect 72 -373 76 -372
rect 80 -373 84 -372
rect 88 -373 92 -372
rect 96 -373 100 -372
rect 104 -373 108 -372
rect 112 -373 116 -372
rect 120 -373 124 -372
rect 128 -373 132 -372
rect 136 -373 140 -372
rect 144 -373 148 -372
rect 152 -373 156 -372
rect 160 -373 164 -372
rect 168 -373 172 -372
rect 176 -373 180 -372
rect 184 -373 188 -372
rect 192 -373 196 -372
rect 200 -373 204 -372
rect 209 -372 212 -365
rect 40 -378 44 -377
rect 56 -378 60 -377
rect 72 -378 76 -377
rect 88 -378 92 -377
rect 104 -378 108 -377
rect 120 -378 124 -377
rect 136 -378 140 -377
rect 152 -378 156 -377
rect 168 -378 172 -377
rect 184 -378 188 -377
rect 200 -378 204 -377
rect 216 -380 224 -364
rect 244 -364 247 -348
rect 254 -356 258 -344
rect 261 -356 265 -355
rect 268 -356 272 -344
rect 283 -348 286 -344
rect 287 -351 290 -348
rect 297 -356 301 -344
rect 333 -349 334 -345
rect 341 -353 345 -341
rect 363 -348 373 -345
rect 366 -353 369 -348
rect 386 -353 390 -341
rect 403 -349 404 -345
rect 408 -349 409 -345
rect 418 -348 421 -176
rect 426 -220 429 -160
rect 434 -172 437 -80
rect 442 -172 445 14
rect 450 4 453 14
rect 450 -44 453 0
rect 450 -60 453 -48
rect 450 -76 453 -64
rect 426 -252 429 -224
rect 426 -268 429 -256
rect 426 -284 429 -272
rect 434 -284 437 -176
rect 442 -220 445 -176
rect 450 -204 453 -80
rect 458 -172 461 14
rect 466 -140 469 14
rect 474 -92 477 14
rect 458 -204 461 -176
rect 408 -357 409 -353
rect 254 -372 258 -360
rect 216 -384 220 -380
rect 8 -534 11 -507
rect 19 -398 32 -394
rect 36 -398 48 -394
rect 52 -398 64 -394
rect 68 -398 80 -394
rect 84 -398 96 -394
rect 100 -398 112 -394
rect 116 -398 128 -394
rect 132 -398 144 -394
rect 148 -398 160 -394
rect 164 -398 176 -394
rect 180 -398 192 -394
rect 196 -398 209 -394
rect 15 -556 19 -398
rect 24 -419 27 -415
rect 24 -422 32 -419
rect 40 -419 43 -415
rect 40 -422 48 -419
rect 56 -419 59 -415
rect 56 -422 64 -419
rect 72 -419 75 -415
rect 72 -422 80 -419
rect 88 -419 91 -415
rect 88 -422 96 -419
rect 104 -419 107 -415
rect 104 -422 112 -419
rect 120 -419 123 -415
rect 120 -422 128 -419
rect 136 -419 139 -415
rect 136 -422 144 -419
rect 152 -419 155 -415
rect 152 -422 160 -419
rect 168 -419 171 -415
rect 168 -422 176 -419
rect 184 -419 187 -415
rect 184 -422 192 -419
rect 24 -425 27 -422
rect 40 -425 43 -422
rect 56 -425 59 -422
rect 72 -425 75 -422
rect 88 -425 91 -422
rect 104 -425 107 -422
rect 120 -425 123 -422
rect 136 -425 139 -422
rect 152 -425 155 -422
rect 168 -425 171 -422
rect 184 -425 187 -422
rect 26 -451 32 -447
rect 36 -451 48 -447
rect 52 -451 64 -447
rect 68 -451 80 -447
rect 84 -451 96 -447
rect 100 -451 112 -447
rect 116 -451 128 -447
rect 132 -451 144 -447
rect 148 -451 160 -447
rect 164 -451 176 -447
rect 180 -451 192 -447
rect 216 -447 224 -384
rect 196 -451 224 -447
rect 26 -485 32 -481
rect 40 -459 44 -458
rect 36 -485 48 -481
rect 56 -459 60 -458
rect 52 -485 64 -481
rect 72 -459 76 -458
rect 68 -485 80 -481
rect 88 -459 92 -458
rect 84 -485 96 -481
rect 104 -459 108 -458
rect 100 -485 112 -481
rect 120 -459 124 -458
rect 116 -485 128 -481
rect 136 -459 140 -458
rect 132 -485 144 -481
rect 152 -459 156 -458
rect 148 -485 160 -481
rect 168 -459 172 -458
rect 164 -485 176 -481
rect 184 -459 188 -458
rect 180 -485 192 -481
rect 200 -459 204 -458
rect 216 -481 224 -451
rect 196 -485 220 -481
rect 30 -493 34 -492
rect 38 -493 42 -492
rect 46 -493 50 -492
rect 54 -493 58 -492
rect 62 -493 66 -492
rect 70 -493 74 -492
rect 78 -493 82 -492
rect 86 -493 90 -492
rect 94 -493 98 -492
rect 102 -493 106 -492
rect 110 -493 114 -492
rect 118 -493 122 -492
rect 126 -493 130 -492
rect 134 -493 138 -492
rect 142 -493 146 -492
rect 150 -493 154 -492
rect 158 -493 162 -492
rect 166 -493 170 -492
rect 174 -493 178 -492
rect 182 -493 186 -492
rect 190 -493 194 -492
rect 198 -493 202 -492
rect 38 -498 42 -497
rect 54 -498 58 -497
rect 70 -498 74 -497
rect 86 -498 90 -497
rect 102 -498 106 -497
rect 118 -498 122 -497
rect 134 -498 138 -497
rect 150 -498 154 -497
rect 166 -498 170 -497
rect 182 -498 186 -497
rect 198 -498 202 -497
rect 26 -507 209 -505
rect 23 -508 209 -507
rect 216 -511 224 -485
rect 26 -515 29 -511
rect 33 -515 38 -511
rect 49 -515 54 -511
rect 65 -515 70 -511
rect 81 -515 86 -511
rect 97 -515 102 -511
rect 113 -515 118 -511
rect 129 -515 134 -511
rect 145 -515 150 -511
rect 161 -515 166 -511
rect 177 -515 182 -511
rect 193 -515 198 -511
rect 209 -515 224 -511
rect 38 -522 39 -518
rect 54 -522 55 -518
rect 70 -522 71 -518
rect 86 -522 87 -518
rect 102 -522 103 -518
rect 118 -522 119 -518
rect 134 -522 135 -518
rect 150 -522 151 -518
rect 166 -522 167 -518
rect 182 -522 183 -518
rect 198 -522 199 -518
rect 35 -529 42 -526
rect 51 -529 58 -526
rect 67 -529 74 -526
rect 83 -529 90 -526
rect 99 -529 106 -526
rect 115 -529 122 -526
rect 131 -529 138 -526
rect 147 -529 154 -526
rect 163 -529 170 -526
rect 179 -529 186 -526
rect 195 -529 202 -526
rect 26 -538 209 -536
rect 23 -539 209 -538
rect 216 -542 224 -515
rect 26 -546 29 -542
rect 33 -546 38 -542
rect 49 -546 54 -542
rect 65 -546 70 -542
rect 81 -546 86 -542
rect 97 -546 102 -542
rect 113 -546 118 -542
rect 129 -546 134 -542
rect 145 -546 150 -542
rect 161 -546 166 -542
rect 177 -546 182 -542
rect 193 -546 198 -542
rect 209 -546 224 -542
rect 38 -553 39 -549
rect 54 -553 55 -549
rect 70 -553 71 -549
rect 86 -553 87 -549
rect 102 -553 103 -549
rect 118 -553 119 -549
rect 134 -553 135 -549
rect 150 -553 151 -549
rect 166 -553 167 -549
rect 182 -553 183 -549
rect 198 -553 199 -549
rect 15 -560 29 -556
rect 33 -560 38 -556
rect 49 -560 54 -556
rect 65 -560 70 -556
rect 81 -560 86 -556
rect 97 -560 102 -556
rect 113 -560 118 -556
rect 129 -560 134 -556
rect 145 -560 150 -556
rect 161 -560 166 -556
rect 177 -560 182 -556
rect 193 -560 198 -556
rect 26 -566 209 -563
rect 35 -576 41 -573
rect 51 -576 57 -573
rect 67 -576 73 -573
rect 83 -576 89 -573
rect 99 -576 105 -573
rect 115 -576 121 -573
rect 131 -576 137 -573
rect 147 -576 153 -573
rect 163 -576 169 -573
rect 179 -576 185 -573
rect 195 -576 201 -573
rect 216 -577 224 -546
rect 268 -372 272 -360
rect 228 -563 231 -376
rect 254 -394 258 -376
rect 297 -380 301 -360
rect 341 -380 345 -357
rect 386 -360 390 -357
rect 418 -360 421 -352
rect 426 -360 429 -288
rect 434 -332 437 -288
rect 442 -316 445 -224
rect 442 -332 445 -320
rect 434 -360 437 -336
rect 442 -348 445 -336
rect 442 -360 445 -352
rect 450 -360 453 -208
rect 458 -300 461 -208
rect 458 -360 461 -304
rect 466 -360 469 -144
rect 474 -360 477 -96
rect 482 -188 485 14
rect 490 -92 493 14
rect 498 4 502 6
rect 498 -4 502 0
rect 498 -12 502 -8
rect 498 -20 502 -16
rect 498 -28 502 -24
rect 498 -36 502 -32
rect 498 -44 502 -40
rect 498 -52 502 -48
rect 498 -60 502 -56
rect 498 -68 502 -64
rect 498 -76 502 -72
rect 498 -84 502 -80
rect 498 -92 502 -88
rect 482 -236 485 -192
rect 482 -360 485 -240
rect 490 -360 493 -96
rect 498 -100 502 -96
rect 498 -108 502 -104
rect 498 -116 502 -112
rect 498 -124 502 -120
rect 498 -132 502 -128
rect 498 -140 502 -136
rect 498 -148 502 -144
rect 498 -156 502 -152
rect 498 -164 502 -160
rect 498 -172 502 -168
rect 498 -180 502 -176
rect 498 -188 502 -184
rect 498 -196 502 -192
rect 498 -204 502 -200
rect 498 -212 502 -208
rect 498 -220 502 -216
rect 498 -228 502 -224
rect 498 -236 502 -232
rect 498 -244 502 -240
rect 498 -252 502 -248
rect 498 -260 502 -256
rect 498 -268 502 -264
rect 498 -276 502 -272
rect 498 -284 502 -280
rect 498 -292 502 -288
rect 498 -300 502 -296
rect 498 -308 502 -304
rect 498 -316 502 -312
rect 498 -324 502 -320
rect 498 -332 502 -328
rect 498 -340 502 -336
rect 498 -348 502 -344
rect 498 -356 502 -352
rect 506 -140 509 14
rect 514 -92 517 14
rect 506 -188 509 -144
rect 506 -268 509 -192
rect 506 -360 509 -272
rect 514 -360 517 -96
rect 522 -140 525 14
rect 530 -124 533 14
rect 530 -140 533 -128
rect 522 -360 525 -144
rect 530 -360 533 -144
rect 538 -188 541 14
rect 546 -108 549 14
rect 538 -236 541 -192
rect 538 -268 541 -240
rect 538 -316 541 -272
rect 546 -300 549 -112
rect 538 -360 541 -320
rect 546 -360 549 -304
rect 554 -316 557 14
rect 563 4 567 6
rect 563 -4 567 0
rect 574 -5 575 -1
rect 563 -12 567 -8
rect 574 -13 575 -9
rect 563 -20 567 -16
rect 574 -21 575 -17
rect 563 -28 567 -24
rect 574 -29 575 -25
rect 563 -36 567 -32
rect 574 -37 575 -33
rect 563 -44 567 -40
rect 574 -45 575 -41
rect 563 -52 567 -48
rect 574 -53 575 -49
rect 563 -60 567 -56
rect 574 -61 575 -57
rect 563 -68 567 -64
rect 574 -69 575 -65
rect 563 -76 567 -72
rect 574 -77 575 -73
rect 563 -84 567 -80
rect 574 -85 575 -81
rect 563 -92 567 -88
rect 574 -93 575 -89
rect 563 -100 567 -96
rect 574 -101 575 -97
rect 563 -108 567 -104
rect 574 -109 575 -105
rect 563 -116 567 -112
rect 563 -124 567 -120
rect 563 -132 567 -128
rect 574 -133 575 -129
rect 563 -140 567 -136
rect 574 -141 575 -137
rect 563 -148 567 -144
rect 574 -149 575 -145
rect 563 -156 567 -152
rect 574 -157 575 -153
rect 563 -164 567 -160
rect 574 -165 575 -161
rect 563 -172 567 -168
rect 574 -173 575 -169
rect 563 -180 567 -176
rect 574 -181 575 -177
rect 563 -188 567 -184
rect 574 -189 575 -185
rect 563 -196 567 -192
rect 574 -197 575 -193
rect 563 -204 567 -200
rect 574 -205 575 -201
rect 563 -212 567 -208
rect 574 -213 575 -209
rect 563 -220 567 -216
rect 574 -221 575 -217
rect 563 -228 567 -224
rect 574 -229 575 -225
rect 563 -236 567 -232
rect 574 -237 575 -233
rect 563 -244 567 -240
rect 563 -252 567 -248
rect 563 -260 567 -256
rect 574 -261 575 -257
rect 563 -268 567 -264
rect 574 -269 575 -265
rect 563 -276 567 -272
rect 574 -277 575 -273
rect 563 -284 567 -280
rect 574 -285 575 -281
rect 563 -292 567 -288
rect 574 -293 575 -289
rect 563 -300 567 -296
rect 574 -301 575 -297
rect 563 -308 567 -304
rect 574 -309 575 -305
rect 563 -316 567 -312
rect 574 -317 575 -313
rect 554 -360 557 -320
rect 563 -324 567 -320
rect 574 -325 575 -321
rect 563 -332 567 -328
rect 574 -333 575 -329
rect 563 -340 567 -336
rect 574 -341 575 -337
rect 563 -348 567 -344
rect 574 -349 575 -345
rect 563 -356 567 -352
rect 574 -357 575 -353
rect 386 -364 394 -360
rect 418 -362 422 -360
rect 426 -362 430 -360
rect 434 -362 438 -360
rect 442 -362 446 -360
rect 450 -362 454 -360
rect 458 -362 462 -360
rect 466 -362 470 -360
rect 474 -362 478 -360
rect 482 -362 486 -360
rect 490 -362 494 -360
rect 506 -362 510 -360
rect 514 -362 518 -360
rect 522 -362 526 -360
rect 530 -362 534 -360
rect 538 -362 542 -360
rect 546 -362 550 -360
rect 554 -362 558 -360
rect 379 -386 382 -368
rect 386 -369 394 -368
rect 386 -372 418 -369
rect 390 -373 418 -372
rect 422 -373 434 -369
rect 438 -373 450 -369
rect 454 -373 466 -369
rect 470 -373 482 -369
rect 486 -373 498 -369
rect 502 -373 506 -369
rect 510 -373 522 -369
rect 526 -373 538 -369
rect 542 -373 554 -369
rect 558 -373 570 -369
rect 390 -376 394 -373
rect 236 -535 239 -508
rect 228 -577 231 -567
rect 236 -577 239 -539
rect 371 -577 374 -442
rect 379 -557 382 -390
rect 379 -577 382 -561
rect 386 -573 394 -376
rect 414 -390 422 -387
rect 426 -390 438 -387
rect 442 -390 454 -387
rect 458 -390 470 -387
rect 474 -390 486 -387
rect 490 -390 510 -387
rect 514 -390 526 -387
rect 530 -390 542 -387
rect 546 -390 574 -387
rect 418 -406 421 -403
rect 434 -406 437 -403
rect 450 -406 453 -403
rect 466 -406 469 -403
rect 482 -406 485 -403
rect 506 -406 509 -403
rect 522 -406 525 -403
rect 538 -406 541 -403
rect 418 -413 421 -410
rect 434 -413 437 -410
rect 450 -413 453 -410
rect 466 -413 469 -410
rect 482 -413 485 -410
rect 506 -413 509 -410
rect 522 -413 525 -410
rect 538 -413 541 -410
rect 414 -442 422 -439
rect 426 -442 438 -439
rect 442 -442 454 -439
rect 458 -442 470 -439
rect 474 -442 486 -439
rect 490 -442 510 -439
rect 514 -442 526 -439
rect 530 -442 542 -439
rect 546 -442 558 -439
rect 562 -442 574 -439
rect 410 -471 418 -467
rect 422 -471 434 -467
rect 438 -471 450 -467
rect 454 -471 466 -467
rect 470 -471 482 -467
rect 486 -471 498 -467
rect 502 -471 506 -467
rect 510 -471 522 -467
rect 526 -471 538 -467
rect 542 -471 554 -467
rect 558 -471 570 -467
rect 410 -481 414 -471
rect 430 -478 431 -474
rect 446 -478 447 -474
rect 462 -478 463 -474
rect 478 -478 479 -474
rect 494 -478 495 -474
rect 518 -478 519 -474
rect 534 -478 535 -474
rect 550 -478 551 -474
rect 566 -478 567 -474
rect 414 -485 434 -481
rect 438 -485 450 -481
rect 454 -485 466 -481
rect 470 -485 482 -481
rect 486 -485 498 -481
rect 502 -485 522 -481
rect 526 -485 538 -481
rect 542 -485 554 -481
rect 558 -485 570 -481
rect 418 -536 421 -533
rect 434 -536 437 -533
rect 450 -536 453 -533
rect 466 -536 469 -533
rect 482 -536 485 -533
rect 506 -536 509 -533
rect 522 -536 525 -533
rect 538 -536 541 -533
rect 554 -536 557 -533
rect 418 -543 421 -540
rect 434 -543 437 -540
rect 450 -543 453 -540
rect 466 -543 469 -540
rect 482 -543 485 -540
rect 506 -543 509 -540
rect 522 -543 525 -540
rect 538 -543 541 -540
rect 554 -543 557 -540
rect 414 -560 422 -557
rect 426 -560 438 -557
rect 442 -560 454 -557
rect 458 -560 470 -557
rect 474 -560 486 -557
rect 490 -560 510 -557
rect 514 -560 526 -557
rect 530 -560 542 -557
rect 546 -560 558 -557
rect 562 -560 574 -557
rect 386 -577 418 -573
rect 422 -577 434 -573
rect 438 -577 450 -573
rect 454 -577 466 -573
rect 470 -577 482 -573
rect 486 -577 498 -573
rect 502 -577 506 -573
rect 510 -577 522 -573
rect 526 -577 538 -573
rect 542 -577 554 -573
rect 558 -577 570 -573
<< metal2 >>
rect 8 20 369 23
rect 8 12 11 20
rect 8 -368 11 8
rect 15 -122 19 12
rect 15 -250 19 -126
rect 15 -394 19 -254
rect 23 -114 26 1
rect 23 -242 26 -118
rect 23 -361 26 -246
rect 31 -366 34 12
rect 39 -366 42 12
rect 47 -366 50 12
rect 55 -366 58 12
rect 63 -366 66 12
rect 71 -366 74 12
rect 79 -366 82 12
rect 87 -366 90 12
rect 95 -366 98 12
rect 103 -366 106 12
rect 111 -366 114 12
rect 119 -366 122 12
rect 127 -366 130 12
rect 135 -366 138 12
rect 143 -366 146 12
rect 151 -366 154 12
rect 159 -366 162 12
rect 167 -366 170 12
rect 175 -366 178 12
rect 183 -366 186 12
rect 191 -366 194 12
rect 199 -366 202 12
rect 366 9 369 20
rect 379 22 409 26
rect 379 17 383 22
rect 405 15 565 18
rect 401 9 404 14
rect 366 6 404 9
rect 413 6 498 10
rect 502 6 563 10
rect 233 0 272 3
rect 287 0 304 3
rect 211 -4 225 -3
rect 211 -6 261 -4
rect 222 -7 261 -6
rect 269 -5 272 0
rect 370 -4 404 -1
rect 408 -4 575 -1
rect 269 -8 304 -5
rect 233 -16 272 -13
rect 338 -13 404 -10
rect 408 -12 575 -9
rect 287 -16 304 -13
rect 211 -20 225 -19
rect 211 -22 261 -20
rect 222 -23 261 -22
rect 269 -21 272 -16
rect 370 -20 404 -17
rect 408 -20 575 -17
rect 269 -24 304 -21
rect 233 -32 272 -29
rect 338 -29 404 -26
rect 408 -28 575 -25
rect 287 -32 304 -29
rect 211 -36 225 -35
rect 211 -38 261 -36
rect 222 -39 261 -38
rect 269 -37 272 -32
rect 370 -36 404 -33
rect 408 -36 575 -33
rect 269 -40 304 -37
rect 233 -48 272 -45
rect 338 -45 404 -42
rect 408 -44 575 -41
rect 287 -48 304 -45
rect 211 -52 225 -51
rect 211 -54 261 -52
rect 222 -55 261 -54
rect 269 -53 272 -48
rect 370 -52 404 -49
rect 408 -52 575 -49
rect 269 -56 304 -53
rect 233 -64 272 -61
rect 338 -61 404 -58
rect 408 -60 575 -57
rect 287 -64 304 -61
rect 211 -68 225 -67
rect 211 -70 261 -68
rect 222 -71 261 -70
rect 269 -69 272 -64
rect 370 -68 404 -65
rect 408 -68 575 -65
rect 269 -72 304 -69
rect 233 -80 272 -77
rect 338 -77 404 -74
rect 408 -76 575 -73
rect 287 -80 304 -77
rect 211 -84 225 -83
rect 211 -86 261 -84
rect 222 -87 261 -86
rect 269 -85 272 -80
rect 370 -84 404 -81
rect 408 -84 575 -81
rect 269 -88 304 -85
rect 233 -96 272 -93
rect 338 -93 404 -90
rect 408 -92 575 -89
rect 287 -96 304 -93
rect 211 -100 225 -99
rect 211 -102 261 -100
rect 222 -103 261 -102
rect 269 -101 272 -96
rect 370 -100 404 -97
rect 408 -100 575 -97
rect 269 -104 304 -101
rect 338 -109 404 -106
rect 408 -108 575 -105
rect 390 -120 498 -116
rect 502 -120 563 -116
rect 233 -128 272 -125
rect 287 -128 304 -125
rect 211 -132 225 -131
rect 211 -134 261 -132
rect 222 -135 261 -134
rect 269 -133 272 -128
rect 370 -132 404 -129
rect 408 -132 575 -129
rect 269 -136 304 -133
rect 233 -144 272 -141
rect 338 -141 404 -138
rect 408 -140 575 -137
rect 287 -144 304 -141
rect 211 -148 225 -147
rect 211 -150 261 -148
rect 222 -151 261 -150
rect 269 -149 272 -144
rect 370 -148 404 -145
rect 408 -148 575 -145
rect 269 -152 304 -149
rect 233 -160 272 -157
rect 338 -157 404 -154
rect 408 -156 575 -153
rect 287 -160 304 -157
rect 211 -164 225 -163
rect 211 -166 261 -164
rect 222 -167 261 -166
rect 269 -165 272 -160
rect 370 -164 404 -161
rect 408 -164 575 -161
rect 269 -168 304 -165
rect 233 -176 272 -173
rect 338 -173 404 -170
rect 408 -172 575 -169
rect 287 -176 304 -173
rect 211 -180 225 -179
rect 211 -182 261 -180
rect 222 -183 261 -182
rect 269 -181 272 -176
rect 370 -180 404 -177
rect 408 -180 575 -177
rect 269 -184 304 -181
rect 233 -192 272 -189
rect 338 -189 404 -186
rect 408 -188 575 -185
rect 287 -192 304 -189
rect 211 -196 225 -195
rect 211 -198 261 -196
rect 222 -199 261 -198
rect 269 -197 272 -192
rect 370 -196 404 -193
rect 408 -196 575 -193
rect 269 -200 304 -197
rect 233 -208 272 -205
rect 338 -205 404 -202
rect 408 -204 575 -201
rect 287 -208 304 -205
rect 211 -212 225 -211
rect 211 -214 261 -212
rect 222 -215 261 -214
rect 269 -213 272 -208
rect 370 -212 404 -209
rect 408 -212 575 -209
rect 269 -216 304 -213
rect 233 -224 272 -221
rect 338 -221 404 -218
rect 408 -220 575 -217
rect 287 -224 304 -221
rect 211 -228 225 -227
rect 211 -230 261 -228
rect 222 -231 261 -230
rect 269 -229 272 -224
rect 370 -228 404 -225
rect 408 -228 575 -225
rect 269 -232 304 -229
rect 338 -237 404 -234
rect 408 -236 575 -233
rect 390 -248 498 -244
rect 502 -248 563 -244
rect 233 -256 272 -253
rect 287 -256 304 -253
rect 211 -260 225 -259
rect 211 -262 261 -260
rect 222 -263 261 -262
rect 269 -261 272 -256
rect 370 -260 404 -257
rect 408 -260 575 -257
rect 269 -264 304 -261
rect 233 -272 272 -269
rect 338 -269 404 -266
rect 408 -268 575 -265
rect 287 -272 304 -269
rect 211 -276 225 -275
rect 211 -278 261 -276
rect 222 -279 261 -278
rect 269 -277 272 -272
rect 370 -276 404 -273
rect 408 -276 575 -273
rect 269 -280 304 -277
rect 233 -288 272 -285
rect 338 -285 404 -282
rect 408 -284 575 -281
rect 287 -288 304 -285
rect 211 -292 225 -291
rect 211 -294 261 -292
rect 222 -295 261 -294
rect 269 -293 272 -288
rect 370 -292 404 -289
rect 408 -292 575 -289
rect 269 -296 304 -293
rect 233 -304 272 -301
rect 338 -301 404 -298
rect 408 -300 575 -297
rect 287 -304 304 -301
rect 211 -308 225 -307
rect 211 -310 261 -308
rect 222 -311 261 -310
rect 269 -309 272 -304
rect 370 -308 404 -305
rect 408 -308 575 -305
rect 269 -312 304 -309
rect 233 -320 272 -317
rect 338 -317 404 -314
rect 408 -316 575 -313
rect 287 -320 304 -317
rect 211 -324 225 -323
rect 211 -326 261 -324
rect 222 -327 261 -326
rect 269 -325 272 -320
rect 370 -324 404 -321
rect 408 -324 575 -321
rect 269 -328 304 -325
rect 233 -336 272 -333
rect 338 -333 404 -330
rect 408 -332 575 -329
rect 287 -336 304 -333
rect 211 -340 225 -339
rect 211 -342 261 -340
rect 222 -343 261 -342
rect 269 -341 272 -336
rect 370 -340 404 -337
rect 408 -340 575 -337
rect 269 -344 304 -341
rect 338 -349 404 -346
rect 408 -348 575 -345
rect 287 -352 304 -349
rect 211 -356 225 -355
rect 211 -358 261 -356
rect 222 -359 261 -358
rect 370 -356 404 -353
rect 408 -356 575 -353
rect 31 -369 35 -366
rect 39 -369 43 -366
rect 47 -369 51 -366
rect 55 -369 59 -366
rect 63 -369 67 -366
rect 71 -369 75 -366
rect 79 -369 83 -366
rect 87 -369 91 -366
rect 95 -369 99 -366
rect 103 -369 107 -366
rect 111 -369 115 -366
rect 119 -369 123 -366
rect 127 -369 131 -366
rect 135 -369 139 -366
rect 143 -369 147 -366
rect 151 -369 155 -366
rect 159 -369 163 -366
rect 167 -369 171 -366
rect 175 -369 179 -366
rect 183 -369 187 -366
rect 191 -369 195 -366
rect 199 -369 203 -366
rect 248 -368 379 -365
rect 32 -373 35 -369
rect 40 -373 43 -369
rect 48 -373 51 -369
rect 56 -373 59 -369
rect 64 -373 67 -369
rect 72 -373 75 -369
rect 80 -373 83 -369
rect 88 -373 91 -369
rect 96 -373 99 -369
rect 104 -373 107 -369
rect 112 -373 115 -369
rect 120 -373 123 -369
rect 128 -373 131 -369
rect 136 -373 139 -369
rect 144 -373 147 -369
rect 152 -373 155 -369
rect 160 -373 163 -369
rect 168 -373 171 -369
rect 176 -373 179 -369
rect 184 -373 187 -369
rect 192 -373 195 -369
rect 200 -373 203 -369
rect 213 -376 228 -373
rect 258 -376 268 -372
rect 272 -376 386 -372
rect 32 -418 35 -377
rect 40 -454 43 -377
rect 48 -418 51 -377
rect 56 -454 59 -377
rect 64 -418 67 -377
rect 72 -454 75 -377
rect 80 -418 83 -377
rect 88 -454 91 -377
rect 96 -418 99 -377
rect 104 -454 107 -377
rect 112 -418 115 -377
rect 120 -454 123 -377
rect 128 -418 131 -377
rect 136 -454 139 -377
rect 144 -418 147 -377
rect 152 -454 155 -377
rect 160 -418 163 -377
rect 168 -454 171 -377
rect 176 -418 179 -377
rect 184 -454 187 -377
rect 192 -418 195 -377
rect 200 -454 203 -377
rect 224 -384 297 -380
rect 301 -384 341 -380
rect 383 -390 410 -387
rect 213 -398 254 -394
rect 418 -399 421 -366
rect 434 -399 437 -366
rect 450 -399 453 -366
rect 466 -399 469 -366
rect 482 -399 485 -366
rect 506 -399 509 -366
rect 522 -399 525 -366
rect 538 -399 541 -366
rect 554 -399 557 -366
rect 418 -402 430 -399
rect 434 -402 446 -399
rect 450 -402 462 -399
rect 466 -402 478 -399
rect 482 -402 494 -399
rect 506 -402 518 -399
rect 522 -402 534 -399
rect 538 -402 550 -399
rect 554 -402 566 -399
rect 375 -442 410 -439
rect 40 -476 43 -458
rect 56 -476 59 -458
rect 72 -476 75 -458
rect 88 -476 91 -458
rect 104 -476 107 -458
rect 120 -476 123 -458
rect 136 -476 139 -458
rect 152 -476 155 -458
rect 168 -476 171 -458
rect 184 -476 187 -458
rect 200 -476 203 -458
rect 31 -479 43 -476
rect 47 -479 59 -476
rect 63 -479 75 -476
rect 79 -479 91 -476
rect 95 -479 107 -476
rect 111 -479 123 -476
rect 127 -479 139 -476
rect 143 -479 155 -476
rect 159 -479 171 -476
rect 175 -479 187 -476
rect 191 -479 203 -476
rect 4 -485 22 -481
rect 31 -493 34 -479
rect 47 -493 50 -479
rect 63 -493 66 -479
rect 79 -493 82 -479
rect 95 -493 98 -479
rect 111 -493 114 -479
rect 127 -493 130 -479
rect 143 -493 146 -479
rect 159 -493 162 -479
rect 175 -493 178 -479
rect 191 -493 194 -479
rect 224 -485 410 -481
rect 38 -501 41 -497
rect 54 -501 57 -497
rect 70 -501 73 -497
rect 86 -501 89 -497
rect 102 -501 105 -497
rect 118 -501 121 -497
rect 134 -501 137 -497
rect 150 -501 153 -497
rect 166 -501 169 -497
rect 182 -501 185 -497
rect 198 -501 201 -497
rect 11 -507 22 -504
rect 31 -504 41 -501
rect 47 -504 57 -501
rect 63 -504 73 -501
rect 79 -504 89 -501
rect 95 -504 105 -501
rect 111 -504 121 -501
rect 127 -504 137 -501
rect 143 -504 153 -501
rect 159 -504 169 -501
rect 175 -504 185 -501
rect 191 -504 201 -501
rect 4 -515 22 -511
rect 31 -525 34 -504
rect 11 -538 22 -535
rect 31 -573 34 -529
rect 39 -549 42 -522
rect 47 -525 50 -504
rect 39 -577 42 -553
rect 47 -573 50 -529
rect 55 -549 58 -522
rect 63 -525 66 -504
rect 55 -577 58 -553
rect 63 -573 66 -529
rect 71 -549 74 -522
rect 79 -525 82 -504
rect 71 -577 74 -553
rect 79 -573 82 -529
rect 87 -549 90 -522
rect 95 -525 98 -504
rect 87 -577 90 -553
rect 95 -573 98 -529
rect 103 -549 106 -522
rect 111 -525 114 -504
rect 103 -577 106 -553
rect 111 -573 114 -529
rect 119 -549 122 -522
rect 127 -525 130 -504
rect 119 -577 122 -553
rect 127 -573 130 -529
rect 135 -549 138 -522
rect 143 -525 146 -504
rect 135 -577 138 -553
rect 143 -573 146 -529
rect 151 -549 154 -522
rect 159 -525 162 -504
rect 151 -577 154 -553
rect 159 -573 162 -529
rect 167 -549 170 -522
rect 175 -525 178 -504
rect 167 -577 170 -553
rect 175 -573 178 -529
rect 183 -549 186 -522
rect 191 -525 194 -504
rect 213 -508 235 -505
rect 418 -509 421 -410
rect 427 -474 430 -402
rect 434 -509 437 -410
rect 443 -474 446 -402
rect 450 -509 453 -410
rect 459 -474 462 -402
rect 466 -509 469 -410
rect 475 -474 478 -402
rect 482 -509 485 -410
rect 491 -474 494 -402
rect 506 -509 509 -410
rect 515 -474 518 -402
rect 522 -509 525 -410
rect 531 -474 534 -402
rect 538 -509 541 -410
rect 547 -474 550 -402
rect 563 -474 566 -402
rect 418 -512 429 -509
rect 434 -512 445 -509
rect 450 -512 461 -509
rect 466 -512 477 -509
rect 482 -512 493 -509
rect 506 -512 517 -509
rect 522 -512 533 -509
rect 538 -512 549 -509
rect 183 -577 186 -553
rect 191 -573 194 -529
rect 199 -549 202 -522
rect 213 -539 235 -536
rect 199 -577 202 -553
rect 383 -560 410 -557
rect 213 -566 228 -563
rect 418 -577 421 -540
rect 426 -577 429 -512
rect 434 -577 437 -540
rect 442 -577 445 -512
rect 450 -577 453 -540
rect 458 -577 461 -512
rect 466 -577 469 -540
rect 474 -577 477 -512
rect 482 -577 485 -540
rect 490 -577 493 -512
rect 506 -577 509 -540
rect 514 -577 517 -512
rect 522 -577 525 -540
rect 530 -577 533 -512
rect 538 -577 541 -540
rect 546 -577 549 -512
rect 554 -577 557 -540
<< ntransistor >>
rect 39 -6 41 -2
rect 39 -14 41 -10
rect 55 -14 57 -10
rect 63 -14 65 -10
rect 39 -22 41 -18
rect 47 -22 49 -18
rect 39 -30 41 -26
rect 39 -38 41 -34
rect 39 -46 41 -42
rect 39 -54 41 -50
rect 39 -62 41 -58
rect 39 -70 41 -66
rect 39 -78 41 -74
rect 39 -86 41 -82
rect 39 -158 41 -154
rect 55 -38 57 -34
rect 39 -166 41 -162
rect 47 -166 49 -162
rect 39 -174 41 -170
rect 39 -206 41 -202
rect 39 -222 41 -218
rect 39 -230 41 -226
rect 39 -262 41 -258
rect 39 -278 41 -274
rect 39 -286 41 -282
rect 39 -294 41 -290
rect 39 -326 41 -322
rect 39 -334 41 -330
rect 39 -342 41 -338
rect 39 -350 41 -346
rect 39 -358 41 -354
rect 71 -22 73 -18
rect 63 -158 65 -154
rect 79 -30 81 -26
rect 103 -6 105 -2
rect 111 -6 113 -2
rect 95 -54 97 -50
rect 87 -62 89 -58
rect 87 -78 89 -74
rect 127 -6 129 -2
rect 135 -14 137 -10
rect 135 -22 137 -18
rect 151 -6 153 -2
rect 151 -14 153 -10
rect 151 -30 153 -26
rect 135 -38 137 -34
rect 143 -38 145 -34
rect 119 -46 121 -42
rect 127 -46 129 -42
rect 127 -54 129 -50
rect 127 -62 129 -58
rect 151 -46 153 -42
rect 151 -54 153 -50
rect 167 -6 169 -2
rect 167 -14 169 -10
rect 167 -22 169 -18
rect 183 -6 185 -2
rect 183 -14 185 -10
rect 167 -30 169 -26
rect 175 -30 177 -26
rect 167 -38 169 -34
rect 167 -46 169 -42
rect 167 -54 169 -50
rect 151 -62 153 -58
rect 159 -62 161 -58
rect 135 -70 137 -66
rect 143 -70 145 -66
rect 127 -78 129 -74
rect 127 -86 129 -82
rect 127 -94 129 -90
rect 159 -70 161 -66
rect 151 -78 153 -74
rect 236 5 240 7
rect 276 5 280 7
rect 199 -6 201 -2
rect 247 -3 251 -1
rect 373 0 383 2
rect 268 -3 272 -1
rect 199 -14 201 -10
rect 236 -11 240 -9
rect 418 -3 422 -1
rect 450 -3 454 -1
rect 393 -8 403 -6
rect 276 -11 280 -9
rect 199 -22 201 -18
rect 247 -19 251 -17
rect 418 -11 422 -9
rect 426 -11 430 -9
rect 434 -11 438 -9
rect 373 -16 383 -14
rect 268 -19 272 -17
rect 191 -30 193 -26
rect 183 -38 185 -34
rect 183 -62 185 -58
rect 175 -70 177 -66
rect 167 -78 169 -74
rect 175 -78 177 -74
rect 151 -86 153 -82
rect 159 -86 161 -82
rect 151 -94 153 -90
rect 159 -94 161 -90
rect 135 -102 137 -98
rect 143 -102 145 -98
rect 135 -110 137 -106
rect 143 -110 145 -106
rect 135 -134 137 -130
rect 143 -134 145 -130
rect 127 -142 129 -138
rect 127 -150 129 -146
rect 135 -158 137 -154
rect 135 -166 137 -162
rect 127 -174 129 -170
rect 135 -182 137 -178
rect 159 -102 161 -98
rect 159 -110 161 -106
rect 159 -134 161 -130
rect 151 -142 153 -138
rect 151 -150 153 -146
rect 236 -27 240 -25
rect 418 -19 422 -17
rect 393 -24 403 -22
rect 276 -27 280 -25
rect 247 -35 251 -33
rect 434 -27 438 -25
rect 373 -32 383 -30
rect 268 -35 272 -33
rect 199 -46 201 -42
rect 236 -43 240 -41
rect 418 -35 422 -33
rect 393 -40 403 -38
rect 276 -43 280 -41
rect 199 -54 201 -50
rect 247 -51 251 -49
rect 426 -43 430 -41
rect 450 -43 454 -41
rect 373 -48 383 -46
rect 268 -51 272 -49
rect 191 -70 193 -66
rect 183 -86 185 -82
rect 236 -59 240 -57
rect 426 -51 430 -49
rect 450 -51 454 -49
rect 393 -56 403 -54
rect 276 -59 280 -57
rect 247 -67 251 -65
rect 418 -59 422 -57
rect 434 -59 438 -57
rect 450 -59 454 -57
rect 373 -64 383 -62
rect 268 -67 272 -65
rect 236 -75 240 -73
rect 450 -67 454 -65
rect 393 -72 403 -70
rect 276 -75 280 -73
rect 199 -86 201 -82
rect 247 -83 251 -81
rect 418 -75 422 -73
rect 426 -75 430 -73
rect 373 -80 383 -78
rect 268 -83 272 -81
rect 183 -94 185 -90
rect 191 -94 193 -90
rect 183 -102 185 -98
rect 191 -102 193 -98
rect 175 -110 177 -106
rect 175 -134 177 -130
rect 167 -142 169 -138
rect 175 -142 177 -138
rect 167 -150 169 -146
rect 159 -158 161 -154
rect 151 -174 153 -170
rect 167 -174 169 -170
rect 151 -182 153 -178
rect 159 -182 161 -178
rect 135 -190 137 -186
rect 143 -190 145 -186
rect 135 -198 137 -194
rect 143 -198 145 -194
rect 127 -206 129 -202
rect 135 -214 137 -210
rect 151 -206 153 -202
rect 151 -214 153 -210
rect 135 -222 137 -218
rect 143 -222 145 -218
rect 135 -230 137 -226
rect 135 -238 137 -234
rect 135 -270 137 -266
rect 135 -286 137 -282
rect 135 -294 137 -290
rect 191 -110 193 -106
rect 236 -91 240 -89
rect 434 -83 438 -81
rect 450 -83 454 -81
rect 393 -88 403 -86
rect 276 -91 280 -89
rect 247 -99 251 -97
rect 474 -91 478 -89
rect 490 -91 494 -89
rect 373 -96 383 -94
rect 268 -99 272 -97
rect 514 -99 518 -97
rect 393 -104 403 -102
rect 546 -107 550 -105
rect 236 -123 240 -121
rect 276 -123 280 -121
rect 199 -134 201 -130
rect 247 -131 251 -129
rect 373 -128 383 -126
rect 268 -131 272 -129
rect 191 -142 193 -138
rect 183 -150 185 -146
rect 191 -150 193 -146
rect 236 -139 240 -137
rect 530 -131 534 -129
rect 393 -136 403 -134
rect 276 -139 280 -137
rect 247 -147 251 -145
rect 466 -139 470 -137
rect 522 -139 526 -137
rect 373 -144 383 -142
rect 268 -147 272 -145
rect 199 -158 201 -154
rect 236 -155 240 -153
rect 183 -166 185 -162
rect 191 -166 193 -162
rect 183 -174 185 -170
rect 191 -174 193 -170
rect 175 -182 177 -178
rect 167 -190 169 -186
rect 175 -190 177 -186
rect 167 -198 169 -194
rect 175 -198 177 -194
rect 167 -206 169 -202
rect 175 -206 177 -202
rect 167 -214 169 -210
rect 175 -214 177 -210
rect 151 -230 153 -226
rect 159 -230 161 -226
rect 151 -238 153 -234
rect 151 -262 153 -258
rect 151 -270 153 -266
rect 151 -278 153 -274
rect 135 -302 137 -298
rect 143 -302 145 -298
rect 127 -310 129 -306
rect 135 -318 137 -314
rect 175 -222 177 -218
rect 175 -230 177 -226
rect 167 -238 169 -234
rect 167 -262 169 -258
rect 506 -147 510 -145
rect 530 -147 534 -145
rect 393 -152 403 -150
rect 276 -155 280 -153
rect 247 -163 251 -161
rect 418 -155 422 -153
rect 373 -160 383 -158
rect 268 -163 272 -161
rect 236 -171 240 -169
rect 426 -163 430 -161
rect 393 -168 403 -166
rect 276 -171 280 -169
rect 199 -182 201 -178
rect 247 -179 251 -177
rect 418 -171 422 -169
rect 434 -171 438 -169
rect 442 -171 446 -169
rect 373 -176 383 -174
rect 268 -179 272 -177
rect 199 -190 201 -186
rect 236 -187 240 -185
rect 191 -198 193 -194
rect 191 -214 193 -210
rect 458 -179 462 -177
rect 393 -184 403 -182
rect 276 -187 280 -185
rect 247 -195 251 -193
rect 482 -187 486 -185
rect 538 -187 542 -185
rect 373 -192 383 -190
rect 268 -195 272 -193
rect 236 -203 240 -201
rect 506 -195 510 -193
rect 538 -195 542 -193
rect 393 -200 403 -198
rect 276 -203 280 -201
rect 247 -211 251 -209
rect 450 -203 454 -201
rect 373 -208 383 -206
rect 268 -211 272 -209
rect 199 -222 201 -218
rect 236 -219 240 -217
rect 183 -238 185 -234
rect 191 -238 193 -234
rect 183 -262 185 -258
rect 191 -262 193 -258
rect 167 -270 169 -266
rect 175 -270 177 -266
rect 167 -278 169 -274
rect 175 -278 177 -274
rect 159 -286 161 -282
rect 151 -310 153 -306
rect 458 -211 462 -209
rect 393 -216 403 -214
rect 276 -219 280 -217
rect 247 -227 251 -225
rect 426 -219 430 -217
rect 373 -224 383 -222
rect 268 -227 272 -225
rect 442 -227 446 -225
rect 393 -232 403 -230
rect 482 -235 486 -233
rect 538 -235 542 -233
rect 236 -251 240 -249
rect 276 -251 280 -249
rect 247 -259 251 -257
rect 373 -256 383 -254
rect 268 -259 272 -257
rect 199 -270 201 -266
rect 236 -267 240 -265
rect 426 -259 430 -257
rect 393 -264 403 -262
rect 276 -267 280 -265
rect 199 -278 201 -274
rect 247 -275 251 -273
rect 506 -267 510 -265
rect 538 -267 542 -265
rect 373 -272 383 -270
rect 268 -275 272 -273
rect 183 -286 185 -282
rect 191 -286 193 -282
rect 167 -294 169 -290
rect 175 -294 177 -290
rect 167 -310 169 -306
rect 151 -318 153 -314
rect 159 -318 161 -314
rect 135 -326 137 -322
rect 143 -326 145 -322
rect 135 -334 137 -330
rect 135 -342 137 -338
rect 143 -342 145 -338
rect 135 -350 137 -346
rect 135 -358 137 -354
rect 143 -358 145 -354
rect 159 -334 161 -330
rect 167 -342 169 -338
rect 191 -294 193 -290
rect 183 -302 185 -298
rect 183 -310 185 -306
rect 236 -283 240 -281
rect 426 -275 430 -273
rect 393 -280 403 -278
rect 276 -283 280 -281
rect 247 -291 251 -289
rect 426 -283 430 -281
rect 434 -283 438 -281
rect 373 -288 383 -286
rect 268 -291 272 -289
rect 199 -302 201 -298
rect 236 -299 240 -297
rect 191 -318 193 -314
rect 183 -326 185 -322
rect 175 -350 177 -346
rect 434 -291 438 -289
rect 393 -296 403 -294
rect 276 -299 280 -297
rect 247 -307 251 -305
rect 458 -299 462 -297
rect 373 -304 383 -302
rect 268 -307 272 -305
rect 236 -315 240 -313
rect 546 -307 550 -305
rect 393 -312 403 -310
rect 276 -315 280 -313
rect 247 -323 251 -321
rect 538 -315 542 -313
rect 554 -315 558 -313
rect 373 -320 383 -318
rect 268 -323 272 -321
rect 199 -334 201 -330
rect 236 -331 240 -329
rect 442 -323 446 -321
rect 393 -328 403 -326
rect 276 -331 280 -329
rect 247 -339 251 -337
rect 434 -331 438 -329
rect 373 -336 383 -334
rect 268 -339 272 -337
rect 199 -350 201 -346
rect 442 -339 446 -337
rect 393 -344 403 -342
rect 276 -347 280 -345
rect 199 -358 201 -354
rect 418 -347 422 -345
rect 373 -352 383 -350
rect 268 -355 272 -353
rect 418 -355 422 -353
rect 442 -355 446 -353
rect 37 -391 39 -378
rect 29 -415 31 -401
rect 53 -391 55 -378
rect 45 -415 47 -401
rect 69 -391 71 -378
rect 61 -415 63 -401
rect 85 -391 87 -378
rect 77 -415 79 -401
rect 101 -391 103 -378
rect 93 -415 95 -401
rect 117 -391 119 -378
rect 109 -415 111 -401
rect 133 -391 135 -378
rect 125 -415 127 -401
rect 149 -391 151 -378
rect 141 -415 143 -401
rect 165 -391 167 -378
rect 157 -415 159 -401
rect 181 -391 183 -378
rect 173 -415 175 -401
rect 197 -391 199 -378
rect 431 -388 433 -376
rect 189 -415 191 -401
rect 423 -403 425 -391
rect 447 -388 449 -376
rect 439 -403 441 -391
rect 463 -388 465 -376
rect 455 -403 457 -391
rect 423 -555 425 -543
rect 479 -388 481 -376
rect 471 -403 473 -391
rect 439 -555 441 -543
rect 38 -563 42 -561
rect 54 -563 58 -561
rect 70 -563 74 -561
rect 86 -563 90 -561
rect 102 -563 106 -561
rect 118 -563 122 -561
rect 134 -563 138 -561
rect 150 -563 154 -561
rect 166 -563 170 -561
rect 182 -563 186 -561
rect 198 -563 202 -561
rect 38 -568 42 -566
rect 54 -568 58 -566
rect 70 -568 74 -566
rect 86 -568 90 -566
rect 102 -568 106 -566
rect 118 -568 122 -566
rect 134 -568 138 -566
rect 150 -568 154 -566
rect 166 -568 170 -566
rect 182 -568 186 -566
rect 198 -568 202 -566
rect 431 -570 433 -558
rect 495 -388 497 -376
rect 487 -403 489 -391
rect 455 -555 457 -543
rect 447 -570 449 -558
rect 519 -388 521 -376
rect 511 -403 513 -391
rect 471 -555 473 -543
rect 463 -570 465 -558
rect 535 -388 537 -376
rect 527 -403 529 -391
rect 487 -555 489 -543
rect 479 -570 481 -558
rect 551 -388 553 -376
rect 543 -403 545 -391
rect 511 -555 513 -543
rect 495 -570 497 -558
rect 527 -555 529 -543
rect 519 -570 521 -558
rect 543 -555 545 -543
rect 535 -570 537 -558
rect 559 -555 561 -543
rect 551 -570 553 -558
rect 567 -570 569 -558
<< ptransistor >>
rect 418 19 422 21
rect 426 19 430 21
rect 434 19 438 21
rect 442 19 446 21
rect 450 19 454 21
rect 458 19 462 21
rect 466 19 470 21
rect 474 19 478 21
rect 482 19 486 21
rect 490 19 494 21
rect 506 19 510 21
rect 514 19 518 21
rect 522 19 526 21
rect 530 19 534 21
rect 538 19 542 21
rect 546 19 550 21
rect 554 19 558 21
rect 9 -6 11 -2
rect 9 -14 11 -10
rect 9 -22 11 -18
rect 9 -30 11 -26
rect 9 -38 11 -34
rect 9 -46 11 -42
rect 9 -54 11 -50
rect 9 -62 11 -58
rect 9 -70 11 -66
rect 9 -78 11 -74
rect 9 -86 11 -82
rect 9 -94 11 -90
rect 9 -102 11 -98
rect 9 -110 11 -106
rect 9 -134 11 -130
rect 9 -142 11 -138
rect 9 -150 11 -146
rect 9 -158 11 -154
rect 9 -166 11 -162
rect 9 -174 11 -170
rect 9 -182 11 -178
rect 9 -190 11 -186
rect 9 -198 11 -194
rect 9 -206 11 -202
rect 9 -214 11 -210
rect 9 -222 11 -218
rect 9 -230 11 -226
rect 9 -238 11 -234
rect 9 -262 11 -258
rect 9 -270 11 -266
rect 9 -278 11 -274
rect 9 -286 11 -282
rect 9 -294 11 -290
rect 9 -302 11 -298
rect 9 -310 11 -306
rect 9 -318 11 -314
rect 9 -326 11 -322
rect 9 -334 11 -330
rect 9 -342 11 -338
rect 9 -350 11 -346
rect 9 -358 11 -354
rect 222 5 226 7
rect 290 5 294 7
rect 222 -3 226 -1
rect 343 0 363 2
rect 290 -3 294 -1
rect 222 -11 226 -9
rect 313 -8 333 -6
rect 290 -11 294 -9
rect 222 -19 226 -17
rect 343 -16 363 -14
rect 290 -19 294 -17
rect 222 -27 226 -25
rect 313 -24 333 -22
rect 290 -27 294 -25
rect 222 -35 226 -33
rect 343 -32 363 -30
rect 290 -35 294 -33
rect 222 -43 226 -41
rect 313 -40 333 -38
rect 290 -43 294 -41
rect 222 -51 226 -49
rect 343 -48 363 -46
rect 290 -51 294 -49
rect 222 -59 226 -57
rect 313 -56 333 -54
rect 290 -59 294 -57
rect 222 -67 226 -65
rect 343 -64 363 -62
rect 290 -67 294 -65
rect 222 -75 226 -73
rect 313 -72 333 -70
rect 290 -75 294 -73
rect 222 -83 226 -81
rect 343 -80 363 -78
rect 290 -83 294 -81
rect 222 -91 226 -89
rect 313 -88 333 -86
rect 290 -91 294 -89
rect 222 -99 226 -97
rect 343 -96 363 -94
rect 290 -99 294 -97
rect 313 -104 333 -102
rect 222 -123 226 -121
rect 290 -123 294 -121
rect 222 -131 226 -129
rect 343 -128 363 -126
rect 290 -131 294 -129
rect 222 -139 226 -137
rect 313 -136 333 -134
rect 290 -139 294 -137
rect 222 -147 226 -145
rect 343 -144 363 -142
rect 290 -147 294 -145
rect 222 -155 226 -153
rect 313 -152 333 -150
rect 290 -155 294 -153
rect 222 -163 226 -161
rect 343 -160 363 -158
rect 290 -163 294 -161
rect 222 -171 226 -169
rect 313 -168 333 -166
rect 290 -171 294 -169
rect 222 -179 226 -177
rect 343 -176 363 -174
rect 290 -179 294 -177
rect 222 -187 226 -185
rect 313 -184 333 -182
rect 290 -187 294 -185
rect 222 -195 226 -193
rect 343 -192 363 -190
rect 290 -195 294 -193
rect 222 -203 226 -201
rect 313 -200 333 -198
rect 290 -203 294 -201
rect 222 -211 226 -209
rect 343 -208 363 -206
rect 290 -211 294 -209
rect 222 -219 226 -217
rect 313 -216 333 -214
rect 290 -219 294 -217
rect 222 -227 226 -225
rect 343 -224 363 -222
rect 290 -227 294 -225
rect 313 -232 333 -230
rect 222 -251 226 -249
rect 290 -251 294 -249
rect 222 -259 226 -257
rect 343 -256 363 -254
rect 290 -259 294 -257
rect 222 -267 226 -265
rect 313 -264 333 -262
rect 290 -267 294 -265
rect 222 -275 226 -273
rect 343 -272 363 -270
rect 290 -275 294 -273
rect 222 -283 226 -281
rect 313 -280 333 -278
rect 290 -283 294 -281
rect 222 -291 226 -289
rect 343 -288 363 -286
rect 290 -291 294 -289
rect 222 -299 226 -297
rect 313 -296 333 -294
rect 290 -299 294 -297
rect 222 -307 226 -305
rect 343 -304 363 -302
rect 290 -307 294 -305
rect 222 -315 226 -313
rect 313 -312 333 -310
rect 290 -315 294 -313
rect 222 -323 226 -321
rect 343 -320 363 -318
rect 290 -323 294 -321
rect 222 -331 226 -329
rect 313 -328 333 -326
rect 290 -331 294 -329
rect 222 -339 226 -337
rect 343 -336 363 -334
rect 290 -339 294 -337
rect 313 -344 333 -342
rect 290 -347 294 -345
rect 343 -352 363 -350
rect 290 -355 294 -353
rect 29 -451 31 -425
rect 45 -451 47 -425
rect 37 -487 39 -461
rect 61 -451 63 -425
rect 53 -487 55 -461
rect 77 -451 79 -425
rect 69 -487 71 -461
rect 93 -451 95 -425
rect 85 -487 87 -461
rect 109 -451 111 -425
rect 101 -487 103 -461
rect 125 -451 127 -425
rect 117 -487 119 -461
rect 141 -451 143 -425
rect 133 -487 135 -461
rect 157 -451 159 -425
rect 149 -487 151 -461
rect 173 -451 175 -425
rect 165 -487 167 -461
rect 189 -451 191 -425
rect 181 -487 183 -461
rect 423 -437 425 -413
rect 439 -437 441 -413
rect 197 -487 199 -461
rect 38 -505 42 -503
rect 54 -505 58 -503
rect 70 -505 74 -503
rect 86 -505 90 -503
rect 102 -505 106 -503
rect 118 -505 122 -503
rect 134 -505 138 -503
rect 150 -505 154 -503
rect 166 -505 170 -503
rect 182 -505 186 -503
rect 198 -505 202 -503
rect 38 -510 42 -508
rect 54 -510 58 -508
rect 70 -510 74 -508
rect 86 -510 90 -508
rect 102 -510 106 -508
rect 118 -510 122 -508
rect 134 -510 138 -508
rect 150 -510 154 -508
rect 166 -510 170 -508
rect 182 -510 186 -508
rect 198 -510 202 -508
rect 431 -464 433 -440
rect 455 -437 457 -413
rect 431 -505 433 -481
rect 38 -536 42 -534
rect 54 -536 58 -534
rect 70 -536 74 -534
rect 86 -536 90 -534
rect 102 -536 106 -534
rect 118 -536 122 -534
rect 134 -536 138 -534
rect 150 -536 154 -534
rect 166 -536 170 -534
rect 182 -536 186 -534
rect 423 -533 425 -509
rect 198 -536 202 -534
rect 38 -541 42 -539
rect 54 -541 58 -539
rect 70 -541 74 -539
rect 86 -541 90 -539
rect 102 -541 106 -539
rect 118 -541 122 -539
rect 134 -541 138 -539
rect 150 -541 154 -539
rect 166 -541 170 -539
rect 182 -541 186 -539
rect 198 -541 202 -539
rect 447 -464 449 -440
rect 471 -437 473 -413
rect 447 -505 449 -481
rect 439 -533 441 -509
rect 463 -464 465 -440
rect 487 -437 489 -413
rect 463 -505 465 -481
rect 455 -533 457 -509
rect 479 -464 481 -440
rect 511 -437 513 -413
rect 479 -505 481 -481
rect 471 -533 473 -509
rect 495 -464 497 -440
rect 527 -437 529 -413
rect 495 -505 497 -481
rect 487 -533 489 -509
rect 519 -464 521 -440
rect 543 -437 545 -413
rect 519 -505 521 -481
rect 511 -533 513 -509
rect 535 -464 537 -440
rect 535 -505 537 -481
rect 527 -533 529 -509
rect 551 -464 553 -440
rect 551 -505 553 -481
rect 543 -533 545 -509
rect 567 -505 569 -481
rect 559 -533 561 -509
<< polycontact >>
rect 565 19 569 23
rect 31 8 35 12
rect 39 8 43 12
rect 47 8 51 12
rect 55 8 59 12
rect 63 8 67 12
rect 71 8 75 12
rect 79 8 83 12
rect 87 8 91 12
rect 95 8 99 12
rect 103 8 107 12
rect 111 8 115 12
rect 119 8 123 12
rect 127 8 131 12
rect 135 8 139 12
rect 143 8 147 12
rect 151 8 155 12
rect 159 8 163 12
rect 167 8 171 12
rect 175 8 179 12
rect 183 8 187 12
rect 191 8 195 12
rect 409 15 413 19
rect 199 8 203 12
rect 7 3 11 7
rect 7 -367 11 -363
rect 243 4 247 8
rect 261 -3 265 1
rect 308 -1 312 3
rect 208 -14 212 -10
rect 243 -12 247 -8
rect 409 -5 413 -1
rect 308 -9 312 -5
rect 570 -5 574 -1
rect 261 -19 265 -15
rect 308 -17 312 -13
rect 409 -13 413 -9
rect 570 -13 574 -9
rect 208 -30 212 -26
rect 243 -28 247 -24
rect 409 -21 413 -17
rect 308 -25 312 -21
rect 570 -21 574 -17
rect 261 -35 265 -31
rect 308 -33 312 -29
rect 409 -29 413 -25
rect 570 -29 574 -25
rect 208 -46 212 -42
rect 243 -44 247 -40
rect 409 -37 413 -33
rect 308 -41 312 -37
rect 570 -37 574 -33
rect 261 -51 265 -47
rect 308 -49 312 -45
rect 409 -45 413 -41
rect 208 -62 212 -58
rect 243 -60 247 -56
rect 570 -45 574 -41
rect 409 -53 413 -49
rect 308 -57 312 -53
rect 570 -53 574 -49
rect 261 -67 265 -63
rect 308 -65 312 -61
rect 409 -61 413 -57
rect 570 -61 574 -57
rect 208 -78 212 -74
rect 243 -76 247 -72
rect 409 -69 413 -65
rect 308 -73 312 -69
rect 570 -69 574 -65
rect 261 -83 265 -79
rect 308 -81 312 -77
rect 409 -77 413 -73
rect 208 -94 212 -90
rect 243 -92 247 -88
rect 570 -77 574 -73
rect 409 -85 413 -81
rect 308 -89 312 -85
rect 570 -85 574 -81
rect 261 -99 265 -95
rect 308 -97 312 -93
rect 409 -93 413 -89
rect 570 -93 574 -89
rect 208 -110 212 -106
rect 409 -101 413 -97
rect 308 -105 312 -101
rect 570 -101 574 -97
rect 409 -109 413 -105
rect 570 -109 574 -105
rect 243 -124 247 -120
rect 261 -131 265 -127
rect 308 -129 312 -125
rect 208 -142 212 -138
rect 243 -140 247 -136
rect 409 -133 413 -129
rect 308 -137 312 -133
rect 570 -133 574 -129
rect 261 -147 265 -143
rect 308 -145 312 -141
rect 409 -141 413 -137
rect 570 -141 574 -137
rect 208 -158 212 -154
rect 243 -156 247 -152
rect 409 -149 413 -145
rect 308 -153 312 -149
rect 570 -149 574 -145
rect 261 -163 265 -159
rect 308 -161 312 -157
rect 409 -157 413 -153
rect 570 -157 574 -153
rect 208 -174 212 -170
rect 243 -172 247 -168
rect 409 -165 413 -161
rect 308 -169 312 -165
rect 570 -165 574 -161
rect 261 -179 265 -175
rect 308 -177 312 -173
rect 409 -173 413 -169
rect 570 -173 574 -169
rect 208 -190 212 -186
rect 243 -188 247 -184
rect 409 -181 413 -177
rect 308 -185 312 -181
rect 570 -181 574 -177
rect 261 -195 265 -191
rect 308 -193 312 -189
rect 409 -189 413 -185
rect 208 -206 212 -202
rect 243 -204 247 -200
rect 570 -189 574 -185
rect 409 -197 413 -193
rect 308 -201 312 -197
rect 570 -197 574 -193
rect 261 -211 265 -207
rect 308 -209 312 -205
rect 409 -205 413 -201
rect 570 -205 574 -201
rect 208 -222 212 -218
rect 243 -220 247 -216
rect 409 -213 413 -209
rect 308 -217 312 -213
rect 570 -213 574 -209
rect 261 -227 265 -223
rect 308 -225 312 -221
rect 409 -221 413 -217
rect 570 -221 574 -217
rect 208 -238 212 -234
rect 409 -229 413 -225
rect 308 -233 312 -229
rect 570 -229 574 -225
rect 409 -237 413 -233
rect 570 -237 574 -233
rect 243 -252 247 -248
rect 261 -259 265 -255
rect 308 -257 312 -253
rect 208 -270 212 -266
rect 243 -268 247 -264
rect 409 -261 413 -257
rect 308 -265 312 -261
rect 570 -261 574 -257
rect 261 -275 265 -271
rect 308 -273 312 -269
rect 409 -269 413 -265
rect 570 -269 574 -265
rect 208 -286 212 -282
rect 243 -284 247 -280
rect 409 -277 413 -273
rect 308 -281 312 -277
rect 570 -277 574 -273
rect 261 -291 265 -287
rect 308 -289 312 -285
rect 409 -285 413 -281
rect 570 -285 574 -281
rect 208 -302 212 -298
rect 243 -300 247 -296
rect 409 -293 413 -289
rect 308 -297 312 -293
rect 570 -293 574 -289
rect 261 -307 265 -303
rect 308 -305 312 -301
rect 409 -301 413 -297
rect 570 -301 574 -297
rect 208 -318 212 -314
rect 243 -316 247 -312
rect 409 -309 413 -305
rect 308 -313 312 -309
rect 570 -309 574 -305
rect 261 -323 265 -319
rect 308 -321 312 -317
rect 409 -317 413 -313
rect 570 -317 574 -313
rect 208 -334 212 -330
rect 243 -332 247 -328
rect 409 -325 413 -321
rect 308 -329 312 -325
rect 570 -325 574 -321
rect 261 -339 265 -335
rect 308 -337 312 -333
rect 409 -333 413 -329
rect 570 -333 574 -329
rect 208 -350 212 -346
rect 243 -348 247 -344
rect 409 -341 413 -337
rect 308 -345 312 -341
rect 570 -341 574 -337
rect 261 -355 265 -351
rect 308 -353 312 -349
rect 409 -349 413 -345
rect 570 -349 574 -345
rect 409 -357 413 -353
rect 570 -357 574 -353
rect 426 -366 430 -362
rect 442 -366 446 -362
rect 458 -366 462 -362
rect 474 -366 478 -362
rect 490 -366 494 -362
rect 514 -366 518 -362
rect 530 -366 534 -362
rect 546 -366 550 -362
rect 32 -372 36 -368
rect 40 -372 44 -368
rect 48 -372 52 -368
rect 56 -372 60 -368
rect 64 -372 68 -368
rect 72 -372 76 -368
rect 80 -372 84 -368
rect 88 -372 92 -368
rect 96 -372 100 -368
rect 104 -372 108 -368
rect 112 -372 116 -368
rect 120 -372 124 -368
rect 128 -372 132 -368
rect 136 -372 140 -368
rect 144 -372 148 -368
rect 152 -372 156 -368
rect 160 -372 164 -368
rect 168 -372 172 -368
rect 176 -372 180 -368
rect 184 -372 188 -368
rect 192 -372 196 -368
rect 200 -372 204 -368
rect 422 -390 426 -386
rect 422 -442 426 -438
rect 438 -390 442 -386
rect 30 -492 34 -488
rect 38 -492 42 -488
rect 46 -492 50 -488
rect 54 -492 58 -488
rect 62 -492 66 -488
rect 70 -492 74 -488
rect 78 -492 82 -488
rect 86 -492 90 -488
rect 94 -492 98 -488
rect 102 -492 106 -488
rect 110 -492 114 -488
rect 118 -492 122 -488
rect 126 -492 130 -488
rect 134 -492 138 -488
rect 142 -492 146 -488
rect 150 -492 154 -488
rect 158 -492 162 -488
rect 166 -492 170 -488
rect 174 -492 178 -488
rect 182 -492 186 -488
rect 190 -492 194 -488
rect 198 -492 202 -488
rect 31 -505 35 -501
rect 47 -505 51 -501
rect 63 -505 67 -501
rect 79 -505 83 -501
rect 95 -505 99 -501
rect 111 -505 115 -501
rect 127 -505 131 -501
rect 143 -505 147 -501
rect 159 -505 163 -501
rect 175 -505 179 -501
rect 191 -505 195 -501
rect 438 -442 442 -438
rect 454 -390 458 -386
rect 431 -478 435 -474
rect 34 -522 38 -518
rect 50 -522 54 -518
rect 66 -522 70 -518
rect 82 -522 86 -518
rect 98 -522 102 -518
rect 114 -522 118 -518
rect 130 -522 134 -518
rect 146 -522 150 -518
rect 162 -522 166 -518
rect 178 -522 182 -518
rect 194 -522 198 -518
rect 31 -536 35 -532
rect 47 -536 51 -532
rect 63 -536 67 -532
rect 79 -536 83 -532
rect 95 -536 99 -532
rect 111 -536 115 -532
rect 127 -536 131 -532
rect 143 -536 147 -532
rect 159 -536 163 -532
rect 175 -536 179 -532
rect 191 -536 195 -532
rect 34 -553 38 -549
rect 50 -553 54 -549
rect 66 -553 70 -549
rect 82 -553 86 -549
rect 98 -553 102 -549
rect 114 -553 118 -549
rect 130 -553 134 -549
rect 146 -553 150 -549
rect 162 -553 166 -549
rect 178 -553 182 -549
rect 194 -553 198 -549
rect 422 -560 426 -556
rect 454 -442 458 -438
rect 470 -390 474 -386
rect 447 -478 451 -474
rect 31 -570 35 -566
rect 47 -570 51 -566
rect 63 -570 67 -566
rect 79 -570 83 -566
rect 95 -570 99 -566
rect 111 -570 115 -566
rect 127 -570 131 -566
rect 143 -570 147 -566
rect 159 -570 163 -566
rect 175 -570 179 -566
rect 191 -570 195 -566
rect 438 -560 442 -556
rect 470 -442 474 -438
rect 486 -390 490 -386
rect 463 -478 467 -474
rect 454 -560 458 -556
rect 486 -442 490 -438
rect 510 -390 514 -386
rect 479 -478 483 -474
rect 470 -560 474 -556
rect 510 -442 514 -438
rect 526 -390 530 -386
rect 495 -478 499 -474
rect 486 -560 490 -556
rect 526 -442 530 -438
rect 542 -390 546 -386
rect 519 -478 523 -474
rect 510 -560 514 -556
rect 542 -442 546 -438
rect 535 -478 539 -474
rect 526 -560 530 -556
rect 558 -442 562 -438
rect 551 -478 555 -474
rect 542 -560 546 -556
rect 567 -478 571 -474
rect 558 -560 562 -556
<< ndcontact >>
rect 34 1 38 5
rect 42 -6 46 -2
rect 42 -14 46 -10
rect 50 1 54 5
rect 66 1 70 5
rect 58 -14 62 -10
rect 42 -22 46 -18
rect 42 -30 46 -26
rect 42 -38 46 -34
rect 42 -46 46 -42
rect 42 -54 46 -50
rect 42 -62 46 -58
rect 42 -70 46 -66
rect 42 -78 46 -74
rect 42 -86 46 -82
rect 34 -118 38 -114
rect 42 -158 46 -154
rect 58 -38 62 -34
rect 50 -118 54 -114
rect 42 -166 46 -162
rect 42 -174 46 -170
rect 42 -206 46 -202
rect 42 -222 46 -218
rect 42 -230 46 -226
rect 34 -246 38 -242
rect 42 -262 46 -258
rect 42 -278 46 -274
rect 42 -286 46 -282
rect 42 -294 46 -290
rect 42 -326 46 -322
rect 42 -334 46 -330
rect 42 -342 46 -338
rect 42 -350 46 -346
rect 42 -358 46 -354
rect 34 -365 38 -361
rect 50 -246 54 -242
rect 50 -365 54 -361
rect 74 -22 78 -18
rect 66 -118 70 -114
rect 58 -158 62 -154
rect 66 -246 70 -242
rect 66 -365 70 -361
rect 82 1 86 5
rect 74 -30 78 -26
rect 98 1 102 5
rect 114 1 118 5
rect 106 -6 110 -2
rect 90 -54 94 -50
rect 90 -62 94 -58
rect 90 -78 94 -74
rect 82 -118 86 -114
rect 82 -246 86 -242
rect 82 -365 86 -361
rect 98 -118 102 -114
rect 98 -246 102 -242
rect 98 -365 102 -361
rect 130 1 134 5
rect 122 -6 126 -2
rect 138 -14 142 -10
rect 138 -22 142 -18
rect 146 1 150 5
rect 154 -6 158 -2
rect 154 -14 158 -10
rect 154 -30 158 -26
rect 138 -38 142 -34
rect 122 -46 126 -42
rect 114 -118 118 -114
rect 114 -246 118 -242
rect 114 -365 118 -361
rect 122 -54 126 -50
rect 122 -62 126 -58
rect 154 -46 158 -42
rect 154 -54 158 -50
rect 162 1 166 5
rect 170 -6 174 -2
rect 170 -14 174 -10
rect 170 -22 174 -18
rect 178 1 182 5
rect 186 -6 190 -2
rect 186 -14 190 -10
rect 170 -30 174 -26
rect 170 -38 174 -34
rect 170 -46 174 -42
rect 170 -54 174 -50
rect 154 -62 158 -58
rect 138 -70 142 -66
rect 122 -78 126 -74
rect 122 -86 126 -82
rect 122 -94 126 -90
rect 154 -70 158 -66
rect 154 -78 158 -74
rect 194 1 198 5
rect 236 8 240 12
rect 276 8 280 12
rect 202 -6 206 -2
rect 373 3 383 7
rect 418 0 422 4
rect 202 -14 206 -10
rect 236 -8 240 -4
rect 250 -8 254 -4
rect 268 -8 272 -4
rect 276 -8 280 -4
rect 450 0 454 4
rect 373 -5 386 -1
rect 390 -5 401 -1
rect 498 -8 502 -4
rect 563 -8 567 -4
rect 202 -22 206 -18
rect 373 -13 383 -9
rect 393 -13 403 -9
rect 418 -16 422 -12
rect 426 -16 430 -12
rect 434 -16 438 -12
rect 186 -30 190 -26
rect 186 -38 190 -34
rect 186 -62 190 -58
rect 170 -70 174 -66
rect 170 -78 174 -74
rect 154 -86 158 -82
rect 154 -94 158 -90
rect 138 -102 142 -98
rect 138 -110 142 -106
rect 130 -118 134 -114
rect 146 -118 150 -114
rect 138 -134 142 -130
rect 122 -142 126 -138
rect 122 -150 126 -146
rect 138 -158 142 -154
rect 138 -166 142 -162
rect 122 -174 126 -170
rect 138 -182 142 -178
rect 154 -102 158 -98
rect 154 -110 158 -106
rect 162 -118 166 -114
rect 154 -134 158 -130
rect 154 -142 158 -138
rect 154 -150 158 -146
rect 236 -24 240 -20
rect 250 -24 254 -20
rect 268 -24 272 -20
rect 276 -24 280 -20
rect 373 -21 386 -17
rect 390 -21 401 -17
rect 498 -24 502 -20
rect 563 -24 567 -20
rect 373 -29 383 -25
rect 393 -29 403 -25
rect 418 -32 422 -28
rect 434 -32 438 -28
rect 202 -46 206 -42
rect 236 -40 240 -36
rect 250 -40 254 -36
rect 268 -40 272 -36
rect 276 -40 280 -36
rect 373 -37 386 -33
rect 390 -37 401 -33
rect 498 -40 502 -36
rect 563 -40 567 -36
rect 202 -54 206 -50
rect 373 -45 383 -41
rect 393 -45 403 -41
rect 426 -48 430 -44
rect 186 -70 190 -66
rect 186 -86 190 -82
rect 236 -56 240 -52
rect 250 -56 254 -52
rect 268 -56 272 -52
rect 276 -56 280 -52
rect 450 -48 454 -44
rect 373 -53 386 -49
rect 390 -53 401 -49
rect 498 -56 502 -52
rect 563 -56 567 -52
rect 373 -61 383 -57
rect 393 -61 403 -57
rect 418 -64 422 -60
rect 434 -64 438 -60
rect 450 -64 454 -60
rect 236 -72 240 -68
rect 250 -72 254 -68
rect 268 -72 272 -68
rect 276 -72 280 -68
rect 373 -69 386 -65
rect 390 -69 401 -65
rect 498 -72 502 -68
rect 563 -72 567 -68
rect 202 -86 206 -82
rect 373 -77 383 -73
rect 393 -77 403 -73
rect 418 -80 422 -76
rect 426 -80 430 -76
rect 434 -80 438 -76
rect 186 -94 190 -90
rect 186 -102 190 -98
rect 170 -110 174 -106
rect 178 -118 182 -114
rect 170 -134 174 -130
rect 170 -142 174 -138
rect 170 -150 174 -146
rect 154 -158 158 -154
rect 154 -174 158 -170
rect 170 -174 174 -170
rect 154 -182 158 -178
rect 138 -190 142 -186
rect 138 -198 142 -194
rect 122 -206 126 -202
rect 138 -214 142 -210
rect 154 -206 158 -202
rect 154 -214 158 -210
rect 138 -222 142 -218
rect 138 -230 142 -226
rect 138 -238 142 -234
rect 130 -246 134 -242
rect 138 -270 142 -266
rect 138 -286 142 -282
rect 138 -294 142 -290
rect 186 -110 190 -106
rect 194 -118 198 -114
rect 236 -88 240 -84
rect 250 -88 254 -84
rect 268 -88 272 -84
rect 276 -88 280 -84
rect 450 -80 454 -76
rect 373 -85 386 -81
rect 390 -85 401 -81
rect 498 -88 502 -84
rect 563 -88 567 -84
rect 373 -93 383 -89
rect 393 -93 403 -89
rect 474 -96 478 -92
rect 490 -96 494 -92
rect 514 -96 518 -92
rect 250 -104 254 -100
rect 268 -104 272 -100
rect 373 -101 386 -97
rect 390 -101 401 -97
rect 498 -104 502 -100
rect 563 -104 567 -100
rect 393 -109 403 -105
rect 546 -112 550 -108
rect 236 -120 240 -116
rect 276 -120 280 -116
rect 202 -134 206 -130
rect 373 -125 383 -121
rect 530 -128 534 -124
rect 186 -142 190 -138
rect 186 -150 190 -146
rect 236 -136 240 -132
rect 250 -136 254 -132
rect 268 -136 272 -132
rect 276 -136 280 -132
rect 373 -133 386 -129
rect 390 -133 401 -129
rect 498 -136 502 -132
rect 563 -136 567 -132
rect 373 -141 383 -137
rect 393 -141 403 -137
rect 466 -144 470 -140
rect 506 -144 510 -140
rect 522 -144 526 -140
rect 530 -144 534 -140
rect 202 -158 206 -154
rect 236 -152 240 -148
rect 250 -152 254 -148
rect 268 -152 272 -148
rect 276 -152 280 -148
rect 186 -166 190 -162
rect 186 -174 190 -170
rect 170 -182 174 -178
rect 170 -190 174 -186
rect 170 -198 174 -194
rect 170 -206 174 -202
rect 170 -214 174 -210
rect 154 -230 158 -226
rect 154 -238 158 -234
rect 146 -246 150 -242
rect 154 -262 158 -258
rect 154 -270 158 -266
rect 154 -278 158 -274
rect 138 -302 142 -298
rect 122 -310 126 -306
rect 138 -318 142 -314
rect 170 -222 174 -218
rect 170 -230 174 -226
rect 170 -238 174 -234
rect 162 -246 166 -242
rect 170 -262 174 -258
rect 373 -149 386 -145
rect 390 -149 401 -145
rect 498 -152 502 -148
rect 563 -152 567 -148
rect 373 -157 383 -153
rect 393 -157 403 -153
rect 418 -160 422 -156
rect 426 -160 430 -156
rect 236 -168 240 -164
rect 250 -168 254 -164
rect 268 -168 272 -164
rect 276 -168 280 -164
rect 373 -165 386 -161
rect 390 -165 401 -161
rect 498 -168 502 -164
rect 563 -168 567 -164
rect 202 -182 206 -178
rect 373 -173 383 -169
rect 393 -173 403 -169
rect 418 -176 422 -172
rect 434 -176 438 -172
rect 442 -176 446 -172
rect 458 -176 462 -172
rect 202 -190 206 -186
rect 236 -184 240 -180
rect 250 -184 254 -180
rect 268 -184 272 -180
rect 276 -184 280 -180
rect 186 -198 190 -194
rect 186 -214 190 -210
rect 373 -181 386 -177
rect 390 -181 401 -177
rect 498 -184 502 -180
rect 563 -184 567 -180
rect 373 -189 383 -185
rect 393 -189 403 -185
rect 482 -192 486 -188
rect 506 -192 510 -188
rect 236 -200 240 -196
rect 250 -200 254 -196
rect 268 -200 272 -196
rect 276 -200 280 -196
rect 538 -192 542 -188
rect 373 -197 386 -193
rect 390 -197 401 -193
rect 498 -200 502 -196
rect 563 -200 567 -196
rect 373 -205 383 -201
rect 393 -205 403 -201
rect 450 -208 454 -204
rect 458 -208 462 -204
rect 202 -222 206 -218
rect 236 -216 240 -212
rect 250 -216 254 -212
rect 268 -216 272 -212
rect 276 -216 280 -212
rect 186 -238 190 -234
rect 178 -246 182 -242
rect 194 -246 198 -242
rect 186 -262 190 -258
rect 170 -270 174 -266
rect 170 -278 174 -274
rect 154 -286 158 -282
rect 154 -310 158 -306
rect 373 -213 386 -209
rect 390 -213 401 -209
rect 498 -216 502 -212
rect 563 -216 567 -212
rect 373 -221 383 -217
rect 393 -221 403 -217
rect 426 -224 430 -220
rect 442 -224 446 -220
rect 250 -232 254 -228
rect 268 -232 272 -228
rect 373 -229 386 -225
rect 390 -229 401 -225
rect 498 -232 502 -228
rect 563 -232 567 -228
rect 393 -237 403 -233
rect 482 -240 486 -236
rect 538 -240 542 -236
rect 236 -248 240 -244
rect 276 -248 280 -244
rect 373 -253 383 -249
rect 426 -256 430 -252
rect 202 -270 206 -266
rect 236 -264 240 -260
rect 250 -264 254 -260
rect 268 -264 272 -260
rect 276 -264 280 -260
rect 373 -261 386 -257
rect 390 -261 401 -257
rect 498 -264 502 -260
rect 563 -264 567 -260
rect 202 -278 206 -274
rect 373 -269 383 -265
rect 393 -269 403 -265
rect 426 -272 430 -268
rect 506 -272 510 -268
rect 538 -272 542 -268
rect 186 -286 190 -282
rect 170 -294 174 -290
rect 170 -310 174 -306
rect 154 -318 158 -314
rect 138 -326 142 -322
rect 138 -334 142 -330
rect 138 -342 142 -338
rect 138 -350 142 -346
rect 138 -358 142 -354
rect 130 -365 134 -361
rect 146 -365 150 -361
rect 154 -334 158 -330
rect 170 -342 174 -338
rect 162 -365 166 -361
rect 186 -294 190 -290
rect 186 -302 190 -298
rect 186 -310 190 -306
rect 236 -280 240 -276
rect 250 -280 254 -276
rect 268 -280 272 -276
rect 276 -280 280 -276
rect 373 -277 386 -273
rect 390 -277 401 -273
rect 498 -280 502 -276
rect 563 -280 567 -276
rect 373 -285 383 -281
rect 393 -285 403 -281
rect 426 -288 430 -284
rect 434 -288 438 -284
rect 202 -302 206 -298
rect 236 -296 240 -292
rect 250 -296 254 -292
rect 268 -296 272 -292
rect 276 -296 280 -292
rect 186 -318 190 -314
rect 186 -326 190 -322
rect 170 -350 174 -346
rect 178 -365 182 -361
rect 373 -293 386 -289
rect 390 -293 401 -289
rect 498 -296 502 -292
rect 563 -296 567 -292
rect 373 -301 383 -297
rect 393 -301 403 -297
rect 458 -304 462 -300
rect 546 -304 550 -300
rect 236 -312 240 -308
rect 250 -312 254 -308
rect 268 -312 272 -308
rect 276 -312 280 -308
rect 373 -309 386 -305
rect 390 -309 401 -305
rect 498 -312 502 -308
rect 563 -312 567 -308
rect 373 -317 383 -313
rect 393 -317 403 -313
rect 442 -320 446 -316
rect 538 -320 542 -316
rect 554 -320 558 -316
rect 202 -334 206 -330
rect 236 -328 240 -324
rect 250 -328 254 -324
rect 268 -328 272 -324
rect 276 -328 280 -324
rect 373 -325 386 -321
rect 390 -325 401 -321
rect 498 -328 502 -324
rect 563 -328 567 -324
rect 373 -333 383 -329
rect 393 -333 403 -329
rect 434 -336 438 -332
rect 442 -336 446 -332
rect 202 -350 206 -346
rect 250 -344 254 -340
rect 268 -344 272 -340
rect 276 -344 280 -340
rect 373 -341 386 -337
rect 390 -341 401 -337
rect 498 -344 502 -340
rect 563 -344 567 -340
rect 202 -358 206 -354
rect 373 -349 383 -345
rect 393 -349 403 -345
rect 418 -352 422 -348
rect 194 -365 198 -361
rect 268 -360 272 -356
rect 442 -352 446 -348
rect 373 -357 386 -353
rect 498 -360 502 -356
rect 563 -360 567 -356
rect 32 -394 36 -380
rect 40 -391 44 -378
rect 24 -415 28 -401
rect 32 -415 36 -398
rect 48 -394 52 -380
rect 56 -391 60 -378
rect 40 -415 44 -401
rect 48 -415 52 -398
rect 64 -394 68 -380
rect 72 -391 76 -378
rect 56 -415 60 -401
rect 64 -415 68 -398
rect 80 -394 84 -380
rect 88 -391 92 -378
rect 72 -415 76 -401
rect 80 -415 84 -398
rect 96 -394 100 -380
rect 104 -391 108 -378
rect 88 -415 92 -401
rect 96 -415 100 -398
rect 112 -394 116 -380
rect 120 -391 124 -378
rect 104 -415 108 -401
rect 112 -415 116 -398
rect 128 -394 132 -380
rect 136 -391 140 -378
rect 120 -415 124 -401
rect 128 -415 132 -398
rect 144 -394 148 -380
rect 152 -391 156 -378
rect 136 -415 140 -401
rect 144 -415 148 -398
rect 160 -394 164 -380
rect 168 -391 172 -378
rect 152 -415 156 -401
rect 160 -415 164 -398
rect 176 -394 180 -380
rect 184 -391 188 -378
rect 168 -415 172 -401
rect 176 -415 180 -398
rect 192 -394 196 -380
rect 200 -391 204 -378
rect 434 -383 438 -373
rect 184 -415 188 -401
rect 192 -415 196 -398
rect 418 -403 422 -393
rect 450 -383 454 -373
rect 434 -403 438 -393
rect 466 -383 470 -373
rect 450 -403 454 -393
rect 418 -553 422 -543
rect 38 -560 45 -556
rect 54 -560 61 -556
rect 70 -560 77 -556
rect 86 -560 93 -556
rect 102 -560 109 -556
rect 118 -560 125 -556
rect 134 -560 141 -556
rect 150 -560 157 -556
rect 166 -560 173 -556
rect 182 -560 189 -556
rect 198 -560 205 -556
rect 482 -383 486 -373
rect 466 -403 470 -393
rect 434 -553 438 -543
rect 38 -573 42 -569
rect 54 -573 58 -569
rect 70 -573 74 -569
rect 86 -573 90 -569
rect 102 -573 106 -569
rect 118 -573 122 -569
rect 134 -573 138 -569
rect 150 -573 154 -569
rect 166 -573 170 -569
rect 182 -573 186 -569
rect 198 -573 202 -569
rect 498 -383 502 -373
rect 482 -403 486 -393
rect 450 -553 454 -543
rect 434 -573 438 -563
rect 522 -383 526 -373
rect 506 -403 510 -393
rect 466 -553 470 -543
rect 450 -573 454 -563
rect 538 -383 542 -373
rect 522 -403 526 -393
rect 482 -553 486 -543
rect 466 -573 470 -563
rect 554 -383 558 -373
rect 538 -403 542 -393
rect 506 -553 510 -543
rect 482 -573 486 -563
rect 522 -553 526 -543
rect 498 -573 502 -563
rect 538 -553 542 -543
rect 522 -573 526 -563
rect 554 -553 558 -543
rect 538 -573 542 -563
rect 554 -573 558 -563
rect 570 -573 574 -563
<< pdcontact >>
rect 416 22 560 26
rect 418 14 422 18
rect 426 14 430 18
rect 434 14 438 18
rect 442 14 446 18
rect 450 14 454 18
rect 458 14 462 18
rect 466 14 470 18
rect 474 14 478 18
rect 482 14 486 18
rect 490 14 494 18
rect 506 14 510 18
rect 514 14 518 18
rect 522 14 526 18
rect 530 14 534 18
rect 538 14 542 18
rect 546 14 550 18
rect 554 14 558 18
rect 219 8 226 12
rect 4 -360 8 0
rect 12 -6 16 -2
rect 12 -14 16 -10
rect 12 -22 16 -18
rect 12 -30 16 -26
rect 12 -38 16 -34
rect 12 -46 16 -42
rect 12 -54 16 -50
rect 12 -62 16 -58
rect 12 -70 16 -66
rect 12 -78 16 -74
rect 12 -86 16 -82
rect 12 -94 16 -90
rect 12 -102 16 -98
rect 12 -110 16 -106
rect 12 -134 16 -130
rect 12 -142 16 -138
rect 12 -150 16 -146
rect 12 -158 16 -154
rect 12 -166 16 -162
rect 12 -174 16 -170
rect 12 -182 16 -178
rect 12 -190 16 -186
rect 12 -198 16 -194
rect 12 -206 16 -202
rect 12 -214 16 -210
rect 12 -222 16 -218
rect 12 -230 16 -226
rect 12 -238 16 -234
rect 12 -262 16 -258
rect 12 -270 16 -266
rect 12 -278 16 -274
rect 12 -286 16 -282
rect 12 -294 16 -290
rect 12 -302 16 -298
rect 12 -310 16 -306
rect 12 -318 16 -314
rect 12 -326 16 -322
rect 12 -334 16 -330
rect 12 -342 16 -338
rect 12 -350 16 -346
rect 12 -358 16 -354
rect 222 0 226 4
rect 290 8 297 12
rect 290 0 294 4
rect 348 3 363 7
rect 219 -8 226 -4
rect 222 -16 226 -12
rect 290 -8 297 -4
rect 315 -5 336 -1
rect 340 -5 363 -1
rect 290 -16 294 -12
rect 315 -13 333 -9
rect 348 -13 363 -9
rect 219 -24 226 -20
rect 222 -32 226 -28
rect 290 -24 297 -20
rect 315 -21 336 -17
rect 340 -21 363 -17
rect 290 -32 294 -28
rect 315 -29 333 -25
rect 348 -29 363 -25
rect 219 -40 226 -36
rect 222 -48 226 -44
rect 290 -40 297 -36
rect 315 -37 336 -33
rect 340 -37 363 -33
rect 290 -48 294 -44
rect 315 -45 333 -41
rect 348 -45 363 -41
rect 219 -56 226 -52
rect 222 -64 226 -60
rect 290 -56 297 -52
rect 315 -53 336 -49
rect 340 -53 363 -49
rect 290 -64 294 -60
rect 315 -61 333 -57
rect 348 -61 363 -57
rect 219 -72 226 -68
rect 222 -80 226 -76
rect 290 -72 297 -68
rect 315 -69 336 -65
rect 340 -69 363 -65
rect 290 -80 294 -76
rect 315 -77 333 -73
rect 348 -77 363 -73
rect 219 -88 226 -84
rect 222 -96 226 -92
rect 290 -88 297 -84
rect 315 -85 336 -81
rect 340 -85 363 -81
rect 290 -96 294 -92
rect 315 -93 333 -89
rect 348 -93 363 -89
rect 219 -104 226 -100
rect 290 -104 297 -100
rect 315 -101 336 -97
rect 340 -101 363 -97
rect 315 -109 333 -105
rect 219 -120 226 -116
rect 222 -128 226 -124
rect 290 -120 297 -116
rect 290 -128 294 -124
rect 348 -125 363 -121
rect 219 -136 226 -132
rect 222 -144 226 -140
rect 290 -136 297 -132
rect 315 -133 336 -129
rect 340 -133 363 -129
rect 290 -144 294 -140
rect 315 -141 333 -137
rect 348 -141 363 -137
rect 219 -152 226 -148
rect 222 -160 226 -156
rect 290 -152 297 -148
rect 315 -149 336 -145
rect 340 -149 363 -145
rect 290 -160 294 -156
rect 315 -157 333 -153
rect 348 -157 363 -153
rect 219 -168 226 -164
rect 222 -176 226 -172
rect 290 -168 297 -164
rect 315 -165 336 -161
rect 340 -165 363 -161
rect 290 -176 294 -172
rect 315 -173 333 -169
rect 348 -173 363 -169
rect 219 -184 226 -180
rect 222 -192 226 -188
rect 290 -184 297 -180
rect 315 -181 336 -177
rect 340 -181 363 -177
rect 290 -192 294 -188
rect 315 -189 333 -185
rect 348 -189 363 -185
rect 219 -200 226 -196
rect 222 -208 226 -204
rect 290 -200 297 -196
rect 315 -197 336 -193
rect 340 -197 363 -193
rect 290 -208 294 -204
rect 315 -205 333 -201
rect 348 -205 363 -201
rect 219 -216 226 -212
rect 222 -224 226 -220
rect 290 -216 297 -212
rect 315 -213 336 -209
rect 340 -213 363 -209
rect 290 -224 294 -220
rect 315 -221 333 -217
rect 348 -221 363 -217
rect 219 -232 226 -228
rect 290 -232 297 -228
rect 315 -229 336 -225
rect 340 -229 363 -225
rect 315 -237 333 -233
rect 219 -248 226 -244
rect 222 -256 226 -252
rect 290 -248 297 -244
rect 290 -256 294 -252
rect 348 -253 363 -249
rect 219 -264 226 -260
rect 222 -272 226 -268
rect 290 -264 297 -260
rect 315 -261 336 -257
rect 340 -261 363 -257
rect 290 -272 294 -268
rect 315 -269 333 -265
rect 348 -269 363 -265
rect 219 -280 226 -276
rect 222 -288 226 -284
rect 290 -280 297 -276
rect 315 -277 336 -273
rect 340 -277 363 -273
rect 290 -288 294 -284
rect 315 -285 333 -281
rect 348 -285 363 -281
rect 219 -296 226 -292
rect 222 -304 226 -300
rect 290 -296 297 -292
rect 315 -293 336 -289
rect 340 -293 363 -289
rect 290 -304 294 -300
rect 315 -301 333 -297
rect 348 -301 363 -297
rect 219 -312 226 -308
rect 222 -320 226 -316
rect 290 -312 297 -308
rect 315 -309 336 -305
rect 340 -309 363 -305
rect 290 -320 294 -316
rect 315 -317 333 -313
rect 348 -317 363 -313
rect 219 -328 226 -324
rect 222 -336 226 -332
rect 290 -328 297 -324
rect 315 -325 336 -321
rect 340 -325 363 -321
rect 290 -336 294 -332
rect 315 -333 333 -329
rect 348 -333 363 -329
rect 219 -344 226 -340
rect 290 -344 297 -340
rect 315 -341 336 -337
rect 340 -341 363 -337
rect 290 -352 294 -348
rect 315 -349 333 -345
rect 348 -349 363 -345
rect 290 -360 297 -356
rect 340 -357 363 -353
rect 24 -444 28 -425
rect 32 -454 36 -425
rect 32 -485 36 -458
rect 40 -444 44 -425
rect 40 -478 44 -459
rect 48 -454 52 -425
rect 48 -485 52 -458
rect 56 -444 60 -425
rect 56 -478 60 -459
rect 64 -454 68 -425
rect 64 -485 68 -458
rect 72 -444 76 -425
rect 72 -478 76 -459
rect 80 -454 84 -425
rect 80 -485 84 -458
rect 88 -444 92 -425
rect 88 -478 92 -459
rect 96 -454 100 -425
rect 96 -485 100 -458
rect 104 -444 108 -425
rect 104 -478 108 -459
rect 112 -454 116 -425
rect 112 -485 116 -458
rect 120 -444 124 -425
rect 120 -478 124 -459
rect 128 -454 132 -425
rect 128 -485 132 -458
rect 136 -444 140 -425
rect 136 -478 140 -459
rect 144 -454 148 -425
rect 144 -485 148 -458
rect 152 -444 156 -425
rect 152 -478 156 -459
rect 160 -454 164 -425
rect 160 -485 164 -458
rect 168 -444 172 -425
rect 168 -478 172 -459
rect 176 -454 180 -425
rect 176 -485 180 -458
rect 184 -444 188 -425
rect 184 -478 188 -459
rect 192 -454 196 -425
rect 192 -485 196 -458
rect 418 -435 422 -413
rect 434 -435 438 -413
rect 200 -478 204 -459
rect 38 -502 42 -498
rect 54 -502 58 -498
rect 70 -502 74 -498
rect 86 -502 90 -498
rect 102 -502 106 -498
rect 118 -502 122 -498
rect 134 -502 138 -498
rect 150 -502 154 -498
rect 166 -502 170 -498
rect 182 -502 186 -498
rect 198 -502 202 -498
rect 450 -435 454 -413
rect 434 -467 438 -445
rect 434 -505 438 -481
rect 38 -515 45 -511
rect 54 -515 61 -511
rect 70 -515 77 -511
rect 86 -515 93 -511
rect 102 -515 109 -511
rect 118 -515 125 -511
rect 134 -515 141 -511
rect 150 -515 157 -511
rect 166 -515 173 -511
rect 182 -515 189 -511
rect 198 -515 205 -511
rect 38 -533 42 -529
rect 54 -533 58 -529
rect 70 -533 74 -529
rect 86 -533 90 -529
rect 102 -533 106 -529
rect 118 -533 122 -529
rect 134 -533 138 -529
rect 150 -533 154 -529
rect 166 -533 170 -529
rect 182 -533 186 -529
rect 198 -533 202 -529
rect 418 -533 422 -509
rect 38 -546 45 -542
rect 54 -546 61 -542
rect 70 -546 77 -542
rect 86 -546 93 -542
rect 102 -546 109 -542
rect 118 -546 125 -542
rect 134 -546 141 -542
rect 150 -546 157 -542
rect 166 -546 173 -542
rect 182 -546 189 -542
rect 198 -546 205 -542
rect 466 -435 470 -413
rect 450 -467 454 -445
rect 450 -505 454 -481
rect 434 -533 438 -509
rect 482 -435 486 -413
rect 466 -467 470 -445
rect 466 -505 470 -481
rect 450 -533 454 -509
rect 506 -435 510 -413
rect 482 -467 486 -445
rect 482 -505 486 -481
rect 466 -533 470 -509
rect 522 -435 526 -413
rect 498 -467 502 -445
rect 498 -505 502 -481
rect 482 -533 486 -509
rect 538 -435 542 -413
rect 522 -467 526 -445
rect 522 -505 526 -481
rect 506 -533 510 -509
rect 538 -467 542 -445
rect 538 -505 542 -481
rect 522 -533 526 -509
rect 554 -467 558 -445
rect 554 -505 558 -481
rect 538 -533 542 -509
rect 570 -505 574 -481
rect 554 -533 558 -509
<< m2contact >>
rect 15 12 19 16
rect 31 12 35 16
rect 7 8 11 12
rect 39 12 43 16
rect 47 12 51 16
rect 55 12 59 16
rect 63 12 67 16
rect 71 12 75 16
rect 79 12 83 16
rect 87 12 91 16
rect 95 12 99 16
rect 103 12 107 16
rect 111 12 115 16
rect 119 12 123 16
rect 127 12 131 16
rect 135 12 139 16
rect 143 12 147 16
rect 151 12 155 16
rect 159 12 163 16
rect 167 12 171 16
rect 175 12 179 16
rect 183 12 187 16
rect 191 12 195 16
rect 199 12 203 16
rect 23 1 27 5
rect 207 -6 211 -2
rect 229 0 233 4
rect 261 -8 265 -4
rect 379 13 383 17
rect 283 0 287 4
rect 304 -1 308 3
rect 409 22 413 26
rect 401 14 405 18
rect 565 14 569 18
rect 409 6 413 10
rect 366 -5 370 -1
rect 404 -5 408 -1
rect 207 -22 211 -18
rect 229 -16 233 -12
rect 261 -24 265 -20
rect 283 -16 287 -12
rect 304 -9 308 -5
rect 334 -13 338 -9
rect 304 -17 308 -13
rect 404 -13 408 -9
rect 366 -21 370 -17
rect 404 -21 408 -17
rect 207 -38 211 -34
rect 229 -32 233 -28
rect 261 -40 265 -36
rect 283 -32 287 -28
rect 304 -25 308 -21
rect 334 -29 338 -25
rect 304 -33 308 -29
rect 404 -29 408 -25
rect 366 -37 370 -33
rect 404 -37 408 -33
rect 207 -54 211 -50
rect 229 -48 233 -44
rect 261 -56 265 -52
rect 283 -48 287 -44
rect 304 -41 308 -37
rect 334 -45 338 -41
rect 304 -49 308 -45
rect 404 -45 408 -41
rect 366 -53 370 -49
rect 404 -53 408 -49
rect 207 -70 211 -66
rect 229 -64 233 -60
rect 261 -72 265 -68
rect 283 -64 287 -60
rect 304 -57 308 -53
rect 334 -61 338 -57
rect 304 -65 308 -61
rect 404 -61 408 -57
rect 366 -69 370 -65
rect 404 -69 408 -65
rect 207 -86 211 -82
rect 229 -80 233 -76
rect 261 -88 265 -84
rect 283 -80 287 -76
rect 304 -73 308 -69
rect 334 -77 338 -73
rect 304 -81 308 -77
rect 404 -77 408 -73
rect 366 -85 370 -81
rect 404 -85 408 -81
rect 207 -102 211 -98
rect 229 -96 233 -92
rect 23 -118 27 -114
rect 261 -104 265 -100
rect 283 -96 287 -92
rect 304 -89 308 -85
rect 334 -93 338 -89
rect 304 -97 308 -93
rect 404 -93 408 -89
rect 366 -101 370 -97
rect 404 -101 408 -97
rect 15 -126 19 -122
rect 207 -134 211 -130
rect 229 -128 233 -124
rect 261 -136 265 -132
rect 304 -105 308 -101
rect 334 -109 338 -105
rect 283 -128 287 -124
rect 304 -129 308 -125
rect 404 -109 408 -105
rect 386 -120 390 -116
rect 366 -133 370 -129
rect 404 -133 408 -129
rect 207 -150 211 -146
rect 229 -144 233 -140
rect 261 -152 265 -148
rect 283 -144 287 -140
rect 304 -137 308 -133
rect 334 -141 338 -137
rect 304 -145 308 -141
rect 404 -141 408 -137
rect 366 -149 370 -145
rect 404 -149 408 -145
rect 207 -166 211 -162
rect 229 -160 233 -156
rect 261 -168 265 -164
rect 283 -160 287 -156
rect 304 -153 308 -149
rect 334 -157 338 -153
rect 304 -161 308 -157
rect 404 -157 408 -153
rect 366 -165 370 -161
rect 404 -165 408 -161
rect 207 -182 211 -178
rect 229 -176 233 -172
rect 261 -184 265 -180
rect 283 -176 287 -172
rect 304 -169 308 -165
rect 334 -173 338 -169
rect 304 -177 308 -173
rect 404 -173 408 -169
rect 366 -181 370 -177
rect 404 -181 408 -177
rect 207 -198 211 -194
rect 229 -192 233 -188
rect 261 -200 265 -196
rect 283 -192 287 -188
rect 304 -185 308 -181
rect 334 -189 338 -185
rect 304 -193 308 -189
rect 404 -189 408 -185
rect 366 -197 370 -193
rect 404 -197 408 -193
rect 207 -214 211 -210
rect 229 -208 233 -204
rect 261 -216 265 -212
rect 283 -208 287 -204
rect 304 -201 308 -197
rect 334 -205 338 -201
rect 304 -209 308 -205
rect 404 -205 408 -201
rect 366 -213 370 -209
rect 404 -213 408 -209
rect 207 -230 211 -226
rect 229 -224 233 -220
rect 23 -246 27 -242
rect 261 -232 265 -228
rect 283 -224 287 -220
rect 304 -217 308 -213
rect 334 -221 338 -217
rect 304 -225 308 -221
rect 404 -221 408 -217
rect 366 -229 370 -225
rect 404 -229 408 -225
rect 15 -254 19 -250
rect 207 -262 211 -258
rect 229 -256 233 -252
rect 261 -264 265 -260
rect 304 -233 308 -229
rect 334 -237 338 -233
rect 283 -256 287 -252
rect 304 -257 308 -253
rect 404 -237 408 -233
rect 386 -248 390 -244
rect 366 -261 370 -257
rect 404 -261 408 -257
rect 207 -278 211 -274
rect 229 -272 233 -268
rect 261 -280 265 -276
rect 283 -272 287 -268
rect 304 -265 308 -261
rect 334 -269 338 -265
rect 304 -273 308 -269
rect 404 -269 408 -265
rect 366 -277 370 -273
rect 404 -277 408 -273
rect 207 -294 211 -290
rect 229 -288 233 -284
rect 261 -296 265 -292
rect 283 -288 287 -284
rect 304 -281 308 -277
rect 334 -285 338 -281
rect 304 -289 308 -285
rect 404 -285 408 -281
rect 366 -293 370 -289
rect 404 -293 408 -289
rect 207 -310 211 -306
rect 229 -304 233 -300
rect 261 -312 265 -308
rect 283 -304 287 -300
rect 304 -297 308 -293
rect 334 -301 338 -297
rect 304 -305 308 -301
rect 404 -301 408 -297
rect 366 -309 370 -305
rect 404 -309 408 -305
rect 207 -326 211 -322
rect 229 -320 233 -316
rect 261 -328 265 -324
rect 283 -320 287 -316
rect 304 -313 308 -309
rect 334 -317 338 -313
rect 304 -321 308 -317
rect 404 -317 408 -313
rect 366 -325 370 -321
rect 404 -325 408 -321
rect 207 -342 211 -338
rect 229 -336 233 -332
rect 261 -344 265 -340
rect 283 -336 287 -332
rect 304 -329 308 -325
rect 334 -333 338 -329
rect 304 -337 308 -333
rect 404 -333 408 -329
rect 366 -341 370 -337
rect 404 -341 408 -337
rect 207 -358 211 -354
rect 23 -365 27 -361
rect 7 -372 11 -368
rect 0 -485 4 -481
rect 32 -377 36 -373
rect 40 -377 44 -373
rect 48 -377 52 -373
rect 56 -377 60 -373
rect 64 -377 68 -373
rect 72 -377 76 -373
rect 80 -377 84 -373
rect 88 -377 92 -373
rect 96 -377 100 -373
rect 104 -377 108 -373
rect 112 -377 116 -373
rect 120 -377 124 -373
rect 128 -377 132 -373
rect 136 -377 140 -373
rect 144 -377 148 -373
rect 152 -377 156 -373
rect 160 -377 164 -373
rect 168 -377 172 -373
rect 176 -377 180 -373
rect 184 -377 188 -373
rect 192 -377 196 -373
rect 200 -377 204 -373
rect 209 -376 213 -372
rect 261 -360 265 -356
rect 283 -352 287 -348
rect 304 -345 308 -341
rect 334 -349 338 -345
rect 304 -353 308 -349
rect 404 -349 408 -345
rect 366 -357 370 -353
rect 404 -357 408 -353
rect 244 -368 248 -364
rect 220 -384 224 -380
rect 7 -507 11 -503
rect 0 -515 4 -511
rect 7 -538 11 -534
rect 15 -398 19 -394
rect 209 -398 213 -394
rect 32 -422 36 -418
rect 48 -422 52 -418
rect 64 -422 68 -418
rect 80 -422 84 -418
rect 96 -422 100 -418
rect 112 -422 116 -418
rect 128 -422 132 -418
rect 144 -422 148 -418
rect 160 -422 164 -418
rect 176 -422 180 -418
rect 192 -422 196 -418
rect 22 -485 26 -481
rect 40 -458 44 -454
rect 56 -458 60 -454
rect 72 -458 76 -454
rect 88 -458 92 -454
rect 104 -458 108 -454
rect 120 -458 124 -454
rect 136 -458 140 -454
rect 152 -458 156 -454
rect 168 -458 172 -454
rect 184 -458 188 -454
rect 200 -458 204 -454
rect 220 -485 224 -481
rect 30 -497 34 -493
rect 38 -497 42 -493
rect 46 -497 50 -493
rect 54 -497 58 -493
rect 62 -497 66 -493
rect 70 -497 74 -493
rect 78 -497 82 -493
rect 86 -497 90 -493
rect 94 -497 98 -493
rect 102 -497 106 -493
rect 110 -497 114 -493
rect 118 -497 122 -493
rect 126 -497 130 -493
rect 134 -497 138 -493
rect 142 -497 146 -493
rect 150 -497 154 -493
rect 158 -497 162 -493
rect 166 -497 170 -493
rect 174 -497 178 -493
rect 182 -497 186 -493
rect 190 -497 194 -493
rect 198 -497 202 -493
rect 22 -507 26 -503
rect 209 -508 213 -504
rect 22 -515 26 -511
rect 39 -522 43 -518
rect 55 -522 59 -518
rect 71 -522 75 -518
rect 87 -522 91 -518
rect 103 -522 107 -518
rect 119 -522 123 -518
rect 135 -522 139 -518
rect 151 -522 155 -518
rect 167 -522 171 -518
rect 183 -522 187 -518
rect 199 -522 203 -518
rect 31 -529 35 -525
rect 47 -529 51 -525
rect 63 -529 67 -525
rect 79 -529 83 -525
rect 95 -529 99 -525
rect 111 -529 115 -525
rect 127 -529 131 -525
rect 143 -529 147 -525
rect 159 -529 163 -525
rect 175 -529 179 -525
rect 191 -529 195 -525
rect 22 -538 26 -534
rect 209 -539 213 -535
rect 39 -553 43 -549
rect 55 -553 59 -549
rect 71 -553 75 -549
rect 87 -553 91 -549
rect 103 -553 107 -549
rect 119 -553 123 -549
rect 135 -553 139 -549
rect 151 -553 155 -549
rect 167 -553 171 -549
rect 183 -553 187 -549
rect 199 -553 203 -549
rect 209 -567 213 -563
rect 31 -577 35 -573
rect 47 -577 51 -573
rect 63 -577 67 -573
rect 79 -577 83 -573
rect 95 -577 99 -573
rect 111 -577 115 -573
rect 127 -577 131 -573
rect 143 -577 147 -573
rect 159 -577 163 -573
rect 175 -577 179 -573
rect 191 -577 195 -573
rect 228 -376 232 -372
rect 254 -376 258 -372
rect 268 -376 272 -372
rect 297 -384 301 -380
rect 498 6 502 10
rect 498 -120 502 -116
rect 498 -248 502 -244
rect 563 6 567 10
rect 575 -5 579 -1
rect 575 -13 579 -9
rect 575 -21 579 -17
rect 575 -29 579 -25
rect 575 -37 579 -33
rect 575 -45 579 -41
rect 575 -53 579 -49
rect 575 -61 579 -57
rect 575 -69 579 -65
rect 575 -77 579 -73
rect 575 -85 579 -81
rect 575 -93 579 -89
rect 575 -101 579 -97
rect 575 -109 579 -105
rect 563 -120 567 -116
rect 575 -133 579 -129
rect 575 -141 579 -137
rect 575 -149 579 -145
rect 575 -157 579 -153
rect 575 -165 579 -161
rect 575 -173 579 -169
rect 575 -181 579 -177
rect 575 -189 579 -185
rect 575 -197 579 -193
rect 575 -205 579 -201
rect 575 -213 579 -209
rect 575 -221 579 -217
rect 575 -229 579 -225
rect 575 -237 579 -233
rect 563 -248 567 -244
rect 575 -261 579 -257
rect 575 -269 579 -265
rect 575 -277 579 -273
rect 575 -285 579 -281
rect 575 -293 579 -289
rect 575 -301 579 -297
rect 575 -309 579 -305
rect 575 -317 579 -313
rect 575 -325 579 -321
rect 575 -333 579 -329
rect 575 -341 579 -337
rect 575 -349 579 -345
rect 575 -357 579 -353
rect 341 -384 345 -380
rect 379 -368 383 -364
rect 418 -366 422 -362
rect 434 -366 438 -362
rect 450 -366 454 -362
rect 466 -366 470 -362
rect 482 -366 486 -362
rect 506 -366 510 -362
rect 522 -366 526 -362
rect 538 -366 542 -362
rect 554 -366 558 -362
rect 254 -398 258 -394
rect 386 -376 390 -372
rect 379 -390 383 -386
rect 371 -442 375 -438
rect 235 -508 239 -504
rect 235 -539 239 -535
rect 228 -567 232 -563
rect 379 -561 383 -557
rect 410 -390 414 -386
rect 418 -410 422 -406
rect 434 -410 438 -406
rect 450 -410 454 -406
rect 466 -410 470 -406
rect 482 -410 486 -406
rect 506 -410 510 -406
rect 522 -410 526 -406
rect 538 -410 542 -406
rect 410 -442 414 -438
rect 426 -478 430 -474
rect 442 -478 446 -474
rect 458 -478 462 -474
rect 474 -478 478 -474
rect 490 -478 494 -474
rect 514 -478 518 -474
rect 530 -478 534 -474
rect 546 -478 550 -474
rect 562 -478 566 -474
rect 410 -485 414 -481
rect 418 -540 422 -536
rect 434 -540 438 -536
rect 450 -540 454 -536
rect 466 -540 470 -536
rect 482 -540 486 -536
rect 506 -540 510 -536
rect 522 -540 526 -536
rect 538 -540 542 -536
rect 554 -540 558 -536
rect 410 -561 414 -557
<< psubstratepcontact >>
rect 26 26 206 30
rect 26 -126 30 -122
rect 26 -254 30 -250
rect 42 -126 46 -122
rect 42 -254 46 -250
rect 58 -126 62 -122
rect 58 -254 62 -250
rect 74 -126 78 -122
rect 74 -254 78 -250
rect 90 -126 94 -122
rect 90 -254 94 -250
rect 106 -126 110 -122
rect 106 -254 110 -250
rect 122 -126 126 -122
rect 254 8 258 12
rect 254 -8 258 -4
rect 498 0 502 4
rect 563 0 567 4
rect 386 -5 390 -1
rect 498 -16 502 -12
rect 563 -16 567 -12
rect 138 -126 142 -122
rect 154 -126 158 -122
rect 254 -24 258 -20
rect 386 -21 390 -17
rect 498 -32 502 -28
rect 563 -32 567 -28
rect 254 -40 258 -36
rect 386 -37 390 -33
rect 254 -56 258 -52
rect 498 -48 502 -44
rect 563 -48 567 -44
rect 386 -53 390 -49
rect 498 -64 502 -60
rect 563 -64 567 -60
rect 254 -72 258 -68
rect 386 -69 390 -65
rect 170 -126 174 -122
rect 122 -254 126 -250
rect 138 -254 142 -250
rect 186 -126 190 -122
rect 254 -88 258 -84
rect 498 -80 502 -76
rect 563 -80 567 -76
rect 386 -85 390 -81
rect 498 -96 502 -92
rect 563 -96 567 -92
rect 254 -104 258 -100
rect 386 -101 390 -97
rect 498 -112 502 -108
rect 563 -112 567 -108
rect 254 -120 258 -116
rect 202 -126 206 -122
rect 498 -128 502 -124
rect 563 -128 567 -124
rect 254 -136 258 -132
rect 386 -133 390 -129
rect 498 -144 502 -140
rect 563 -144 567 -140
rect 254 -152 258 -148
rect 154 -254 158 -250
rect 170 -254 174 -250
rect 386 -149 390 -145
rect 498 -160 502 -156
rect 563 -160 567 -156
rect 254 -168 258 -164
rect 386 -165 390 -161
rect 498 -176 502 -172
rect 563 -176 567 -172
rect 254 -184 258 -180
rect 386 -181 390 -177
rect 498 -192 502 -188
rect 254 -200 258 -196
rect 563 -192 567 -188
rect 386 -197 390 -193
rect 498 -208 502 -204
rect 563 -208 567 -204
rect 254 -216 258 -212
rect 186 -254 190 -250
rect 386 -213 390 -209
rect 498 -224 502 -220
rect 563 -224 567 -220
rect 254 -232 258 -228
rect 386 -229 390 -225
rect 498 -240 502 -236
rect 563 -240 567 -236
rect 254 -248 258 -244
rect 202 -254 206 -250
rect 498 -256 502 -252
rect 563 -256 567 -252
rect 254 -264 258 -260
rect 386 -261 390 -257
rect 498 -272 502 -268
rect 563 -272 567 -268
rect 254 -280 258 -276
rect 386 -277 390 -273
rect 498 -288 502 -284
rect 563 -288 567 -284
rect 254 -296 258 -292
rect 386 -293 390 -289
rect 498 -304 502 -300
rect 563 -304 567 -300
rect 254 -312 258 -308
rect 386 -309 390 -305
rect 498 -320 502 -316
rect 563 -320 567 -316
rect 254 -328 258 -324
rect 386 -325 390 -321
rect 498 -336 502 -332
rect 563 -336 567 -332
rect 254 -344 258 -340
rect 386 -341 390 -337
rect 254 -360 258 -356
rect 498 -352 502 -348
rect 563 -352 567 -348
rect 386 -357 390 -353
rect 386 -368 394 -364
rect 418 -373 422 -369
rect 434 -373 438 -369
rect 32 -398 36 -394
rect 48 -398 52 -394
rect 64 -398 68 -394
rect 80 -398 84 -394
rect 96 -398 100 -394
rect 112 -398 116 -394
rect 128 -398 132 -394
rect 144 -398 148 -394
rect 160 -398 164 -394
rect 176 -398 180 -394
rect 450 -373 454 -369
rect 192 -398 196 -394
rect 466 -373 470 -369
rect 482 -373 486 -369
rect 29 -560 33 -556
rect 45 -560 49 -556
rect 61 -560 65 -556
rect 77 -560 81 -556
rect 93 -560 97 -556
rect 109 -560 113 -556
rect 125 -560 129 -556
rect 141 -560 145 -556
rect 157 -560 161 -556
rect 173 -560 177 -556
rect 189 -560 193 -556
rect 205 -560 209 -556
rect 498 -373 502 -369
rect 506 -373 510 -369
rect 522 -373 526 -369
rect 538 -373 542 -369
rect 418 -577 422 -573
rect 434 -577 438 -573
rect 554 -373 558 -369
rect 570 -373 574 -369
rect 450 -577 454 -573
rect 466 -577 470 -573
rect 482 -577 486 -573
rect 498 -577 502 -573
rect 506 -577 510 -573
rect 522 -577 526 -573
rect 538 -577 542 -573
rect 554 -577 558 -573
rect 570 -577 574 -573
<< nsubstratencontact >>
rect 416 26 560 30
rect 215 8 219 12
rect 0 -360 4 0
rect 297 8 301 12
rect 215 -8 219 -4
rect 297 -8 301 -4
rect 336 -5 340 -1
rect 215 -24 219 -20
rect 297 -24 301 -20
rect 336 -21 340 -17
rect 215 -40 219 -36
rect 297 -40 301 -36
rect 336 -37 340 -33
rect 215 -56 219 -52
rect 297 -56 301 -52
rect 336 -53 340 -49
rect 215 -72 219 -68
rect 297 -72 301 -68
rect 336 -69 340 -65
rect 215 -88 219 -84
rect 297 -88 301 -84
rect 336 -85 340 -81
rect 215 -104 219 -100
rect 297 -104 301 -100
rect 336 -101 340 -97
rect 215 -120 219 -116
rect 297 -120 301 -116
rect 215 -136 219 -132
rect 297 -136 301 -132
rect 336 -133 340 -129
rect 215 -152 219 -148
rect 297 -152 301 -148
rect 336 -149 340 -145
rect 215 -168 219 -164
rect 297 -168 301 -164
rect 336 -165 340 -161
rect 215 -184 219 -180
rect 297 -184 301 -180
rect 336 -181 340 -177
rect 215 -200 219 -196
rect 297 -200 301 -196
rect 336 -197 340 -193
rect 215 -216 219 -212
rect 297 -216 301 -212
rect 336 -213 340 -209
rect 215 -232 219 -228
rect 297 -232 301 -228
rect 336 -229 340 -225
rect 215 -248 219 -244
rect 297 -248 301 -244
rect 215 -264 219 -260
rect 297 -264 301 -260
rect 336 -261 340 -257
rect 215 -280 219 -276
rect 297 -280 301 -276
rect 336 -277 340 -273
rect 215 -296 219 -292
rect 297 -296 301 -292
rect 336 -293 340 -289
rect 215 -312 219 -308
rect 297 -312 301 -308
rect 336 -309 340 -305
rect 215 -328 219 -324
rect 297 -328 301 -324
rect 336 -325 340 -321
rect 215 -344 219 -340
rect 297 -344 301 -340
rect 336 -341 340 -337
rect 215 -360 219 -356
rect 297 -360 301 -356
rect 336 -357 340 -353
rect 32 -458 36 -454
rect 48 -458 52 -454
rect 64 -458 68 -454
rect 80 -458 84 -454
rect 96 -458 100 -454
rect 112 -458 116 -454
rect 128 -458 132 -454
rect 144 -458 148 -454
rect 160 -458 164 -454
rect 176 -458 180 -454
rect 192 -458 196 -454
rect 418 -471 422 -467
rect 434 -471 438 -467
rect 29 -515 33 -511
rect 45 -515 49 -511
rect 61 -515 65 -511
rect 77 -515 81 -511
rect 93 -515 97 -511
rect 109 -515 113 -511
rect 125 -515 129 -511
rect 141 -515 145 -511
rect 157 -515 161 -511
rect 173 -515 177 -511
rect 189 -515 193 -511
rect 205 -515 209 -511
rect 29 -546 33 -542
rect 45 -546 49 -542
rect 61 -546 65 -542
rect 77 -546 81 -542
rect 93 -546 97 -542
rect 109 -546 113 -542
rect 125 -546 129 -542
rect 141 -546 145 -542
rect 157 -546 161 -542
rect 173 -546 177 -542
rect 189 -546 193 -542
rect 205 -546 209 -542
rect 450 -471 454 -467
rect 466 -471 470 -467
rect 482 -471 486 -467
rect 498 -471 502 -467
rect 506 -471 510 -467
rect 522 -471 526 -467
rect 538 -471 542 -467
rect 554 -471 558 -467
rect 570 -471 574 -467
<< labels >>
rlabel metal2 40 -555 40 -555 1 RESET
rlabel metal2 56 -555 56 -555 1 req_d
rlabel metal2 72 -555 72 -555 1 req_v
rlabel metal2 88 -555 88 -555 1 ack_out
rlabel metal2 104 -555 104 -555 1 icarry
rlabel metal2 120 -555 120 -555 1 scarry
rlabel metal2 136 -555 136 -555 1 InSt0*
rlabel metal2 152 -555 152 -555 1 InSt1*
rlabel metal2 168 -555 168 -555 1 InSt2*
rlabel metal2 184 -555 184 -555 1 InSt3*
rlabel metal2 200 -555 200 -555 1 InSt4*
rlabel metal1 372 -576 372 -576 1 p1_
rlabel metal1 380 -576 380 -576 1 p1
rlabel metal1 237 -576 237 -576 1 p2_
rlabel metal1 229 -576 229 -576 1 p2
rlabel metal1 390 -576 390 -576 1 GND
rlabel metal1 220 -576 220 -576 1 Vdd
rlabel metal1 419 -535 419 -535 1 OutSt4*
rlabel metal2 427 -535 427 -535 1 OutSt3*
rlabel metal1 435 -535 435 -535 1 OutSt2*
rlabel metal2 443 -535 443 -535 1 OutSt1*
rlabel metal1 451 -535 451 -535 1 OutSt0*
rlabel metal2 459 -535 459 -535 1 ack_in
rlabel metal1 467 -535 467 -535 1 req_Q
rlabel metal2 475 -535 475 -535 1 req_R
rlabel metal1 483 -535 483 -535 1 sreg_reset
rlabel metal2 491 -535 491 -535 1 sreg_rd
rlabel metal1 507 -535 507 -535 1 sreg_wr
rlabel metal2 515 -535 515 -535 1 ireg_reset
rlabel metal1 523 -535 523 -535 1 ireg_rd
rlabel metal2 531 -535 531 -535 1 ireg_wr
rlabel metal1 539 -535 539 -535 1 io_rd
rlabel metal2 547 -535 547 -535 1 reg_rd
rlabel metal1 555 -535 555 -535 1 reg_wr
<< end >>
