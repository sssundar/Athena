magic
tech scmos
timestamp 1434187039
<< polysilicon >>
rect -282 1783 -274 1785
rect -282 1775 -265 1777
rect -214 1774 -199 1776
rect -282 1767 -278 1769
rect -201 1769 -199 1774
rect -282 1759 -280 1767
rect -282 1751 -258 1753
rect -282 1743 -274 1745
rect 132 999 150 1001
rect 132 977 134 999
rect 1227 956 1232 958
rect 1230 946 1232 956
rect 1230 944 1264 946
rect 1288 842 1290 853
rect 1193 694 1264 696
rect 1288 592 1290 603
rect 1193 444 1264 446
rect 1288 342 1290 353
rect 1193 194 1264 196
rect 1288 92 1290 103
rect 1286 57 1329 59
<< metal1 >>
rect -313 1809 -310 1838
rect -277 1809 -274 1830
rect -264 1779 -261 1864
rect -278 1766 -274 1767
rect -258 1755 -255 1847
rect -218 1778 -215 1847
rect -204 1805 -201 1838
rect -173 1805 -170 1830
rect -154 1764 -151 1821
rect -110 1752 -107 1800
rect -110 879 -107 1748
rect -102 1652 -99 1800
rect -110 0 -107 875
rect -102 754 -99 1648
rect -94 1552 -91 1800
rect -102 0 -99 750
rect -94 629 -91 1548
rect -86 1452 -83 1800
rect -94 0 -91 625
rect -86 504 -83 1448
rect -78 1352 -75 1800
rect -86 0 -83 500
rect -78 379 -75 1348
rect -70 1252 -67 1800
rect -78 0 -75 375
rect -70 254 -67 1248
rect -62 1152 -59 1800
rect -70 0 -67 250
rect -62 129 -59 1148
rect -54 1052 -51 1800
rect 1365 1738 1386 1741
rect 1382 1692 1386 1738
rect 1370 1688 1386 1692
rect 1370 1679 1374 1688
rect 1286 1640 1287 1644
rect 1286 1619 1287 1623
rect 1370 1588 1374 1675
rect 1286 1513 1287 1517
rect 1370 1474 1374 1584
rect 1286 1437 1287 1441
rect 1286 1416 1287 1420
rect 1370 1384 1374 1470
rect 1286 1310 1287 1314
rect 1370 1270 1374 1380
rect 1286 1234 1287 1238
rect 1286 1213 1287 1217
rect 1370 1179 1374 1266
rect -62 0 -59 125
rect -54 4 -51 1048
rect 317 1110 327 1113
rect 70 1036 76 1040
rect 102 1036 123 1039
rect 58 988 61 1012
rect 70 994 74 1036
rect 85 1026 88 1033
rect 120 1032 123 1036
rect 120 1029 132 1032
rect 129 994 132 1029
rect 135 1016 138 1036
rect 159 1010 162 1036
rect 142 1007 162 1010
rect 192 1008 196 1036
rect 142 988 145 1007
rect 216 1001 220 1036
rect 154 997 220 1001
rect 317 988 321 1110
rect 1286 1107 1287 1111
rect 1370 1065 1374 1175
rect 1286 1031 1287 1035
rect 1286 1010 1287 1014
rect 1370 974 1374 1061
rect 1223 954 1227 955
rect 1286 904 1287 908
rect 1287 857 1291 858
rect 1370 845 1374 970
rect 1286 806 1287 810
rect 1286 785 1287 789
rect 1370 725 1374 841
rect 1189 690 1193 693
rect 1286 654 1287 658
rect 1287 607 1291 608
rect 1370 594 1374 721
rect 1286 556 1287 560
rect 1286 535 1287 539
rect 1370 475 1374 590
rect 1189 440 1193 443
rect 1286 404 1287 408
rect 1287 357 1291 358
rect 1370 344 1374 471
rect 1286 306 1287 310
rect 1286 285 1287 289
rect 1370 225 1374 340
rect 1189 190 1193 193
rect 1286 154 1287 158
rect 1287 107 1291 108
rect 1333 56 1334 60
rect 1286 35 1287 39
rect 1370 31 1374 221
rect 7 -12 10 0
rect 38 -4 41 8
rect 79 -12 82 0
rect 121 -4 124 8
rect 168 -4 171 8
rect 190 -5 194 0
rect 204 -5 208 1
rect 285 -5 289 0
rect 190 -9 289 -5
rect 317 -4 321 9
rect 204 -12 208 -9
rect 352 -12 355 0
rect 393 -4 397 0
rect 429 -4 432 0
rect 435 -12 438 0
rect 509 -12 513 5
rect 614 -12 617 0
rect 645 -4 648 0
rect 686 -12 689 0
rect 722 -4 725 8
rect 741 -8 744 0
rect 748 -8 751 0
rect 755 -4 758 8
rect 796 -12 799 0
rect 823 -12 826 0
rect 859 -4 862 8
rect 886 -4 889 8
rect 893 -12 896 0
rect 932 -4 935 8
rect 939 -12 942 0
rect 965 -12 968 0
rect 1001 -4 1004 0
rect 1035 -12 1038 0
rect 1071 -4 1074 0
rect 1105 -12 1108 0
rect 1141 -4 1144 0
rect 1175 -12 1178 0
rect 1211 -4 1214 0
rect 1258 -12 1261 0
rect 1294 -4 1297 0
rect 1370 -12 1374 27
rect 1381 1600 1385 1679
rect 1381 1528 1385 1596
rect 1381 1395 1385 1524
rect 1381 1323 1385 1391
rect 1381 1190 1385 1319
rect 1381 1118 1385 1186
rect 1381 985 1385 1114
rect 1381 913 1385 981
rect 1381 765 1385 909
rect 1381 693 1385 761
rect 1381 515 1385 689
rect 1381 443 1385 511
rect 1381 265 1385 439
rect 1381 193 1385 261
rect 1381 91 1385 189
rect 1381 -4 1385 87
<< metal2 >>
rect -313 1880 1367 1884
rect -313 1872 1367 1876
rect -313 1864 -265 1868
rect -261 1864 1367 1868
rect -313 1856 1367 1860
rect -313 1847 -258 1851
rect -254 1847 -218 1851
rect -214 1847 1367 1851
rect -309 1838 -204 1842
rect -200 1838 1367 1842
rect -273 1830 -173 1834
rect -169 1830 1367 1834
rect -313 1821 -155 1825
rect -151 1821 1367 1825
rect -119 1748 -111 1752
rect 1374 1676 1390 1679
rect -119 1648 -103 1652
rect 1287 1644 1390 1646
rect 1291 1642 1390 1644
rect 1287 1618 1291 1619
rect 1287 1615 1390 1618
rect 1385 1596 1390 1600
rect 1374 1585 1390 1588
rect 1275 1573 1393 1577
rect -119 1548 -95 1552
rect 1385 1524 1401 1528
rect 1291 1513 1393 1517
rect 1374 1470 1390 1474
rect -119 1448 -87 1452
rect 1291 1437 1390 1441
rect 1287 1413 1291 1416
rect 1287 1410 1391 1413
rect 1385 1391 1390 1395
rect 1374 1380 1390 1383
rect 1275 1370 1393 1374
rect -119 1348 -79 1352
rect 1385 1319 1390 1323
rect 1291 1310 1393 1314
rect 1374 1266 1390 1269
rect -119 1248 -71 1252
rect 1291 1234 1390 1236
rect 1287 1232 1390 1234
rect 1287 1208 1291 1213
rect 1287 1205 1390 1208
rect 1385 1186 1390 1190
rect 1374 1175 1390 1178
rect 1275 1167 1393 1171
rect -119 1148 -63 1152
rect 1385 1114 1390 1118
rect 1291 1107 1393 1110
rect 1374 1061 1390 1064
rect -119 1048 -55 1052
rect 1287 1027 1393 1031
rect 62 1012 135 1016
rect 72 1004 192 1008
rect 72 988 76 1004
rect 1287 1003 1291 1010
rect 1287 1000 1390 1003
rect 1385 981 1390 985
rect 1374 970 1390 973
rect 1275 964 1393 966
rect 1271 963 1393 964
rect 627 902 631 944
rect 1223 940 1227 950
rect 712 935 979 939
rect 1189 936 1227 940
rect 1385 909 1390 913
rect 991 904 1205 908
rect 365 886 369 901
rect 476 898 704 902
rect 1287 901 1393 904
rect 92 879 96 885
rect 165 882 369 886
rect -106 875 96 879
rect 1189 858 1287 862
rect 627 777 631 819
rect 1189 815 1193 858
rect 1374 841 1390 844
rect 712 810 979 814
rect 1287 810 1390 811
rect 1291 807 1390 810
rect 1287 783 1291 785
rect 991 779 1205 783
rect 1287 780 1390 783
rect 365 761 369 776
rect 476 773 704 777
rect 1385 761 1390 765
rect 92 754 96 760
rect 165 757 369 761
rect -98 750 96 754
rect 1374 721 1390 724
rect 1275 714 1391 717
rect 627 652 631 694
rect 1385 689 1390 693
rect 712 685 979 689
rect 991 654 1205 658
rect 1291 654 1390 658
rect 365 636 369 651
rect 476 648 704 652
rect 92 629 96 635
rect 165 632 369 636
rect -90 625 96 629
rect 1189 608 1287 612
rect 627 527 631 569
rect 1189 565 1193 608
rect 1374 590 1390 594
rect 712 560 979 564
rect 1287 560 1390 561
rect 1291 557 1390 560
rect 1287 533 1291 535
rect 991 529 1205 533
rect 1287 530 1390 533
rect 365 511 369 526
rect 476 523 704 527
rect 1385 511 1391 515
rect 92 504 96 510
rect 165 507 369 511
rect -82 500 96 504
rect 1374 471 1390 474
rect 1275 464 1390 467
rect 627 402 631 444
rect 1385 439 1401 443
rect 712 435 979 439
rect 991 404 1205 408
rect 1291 404 1390 408
rect 365 386 369 401
rect 476 398 704 402
rect 92 379 96 385
rect 165 382 369 386
rect -74 375 96 379
rect 1189 358 1287 362
rect 627 277 631 319
rect 1189 315 1193 358
rect 1374 340 1390 344
rect 712 310 979 314
rect 1287 310 1391 311
rect 1291 307 1391 310
rect 1287 283 1291 285
rect 991 279 1205 283
rect 1287 280 1392 283
rect 365 261 369 276
rect 476 273 704 277
rect 1385 261 1391 265
rect 92 254 96 260
rect 165 257 369 261
rect -66 250 96 254
rect 1374 221 1390 224
rect 1275 214 1390 217
rect 627 152 631 194
rect 1385 189 1401 193
rect 712 185 983 189
rect 991 154 1205 158
rect 1291 154 1390 158
rect 365 136 369 151
rect 476 148 704 152
rect 92 129 96 135
rect 165 132 369 136
rect -58 125 96 129
rect 1189 108 1287 112
rect 1189 65 1193 108
rect 1385 87 1390 91
rect 712 60 983 64
rect 627 27 631 58
rect 1338 56 1390 60
rect 1291 35 1390 39
rect 995 29 1061 33
rect 1065 29 1205 33
rect 1374 27 1390 31
rect 365 11 369 26
rect 476 23 704 27
rect 92 4 96 10
rect 165 7 369 11
rect -50 0 96 4
rect 466 -4 470 0
rect -42 -8 38 -4
rect 42 -8 121 -4
rect 125 -8 168 -4
rect 172 -8 317 -4
rect 321 -8 393 -4
rect 397 -8 428 -4
rect 432 -8 645 -4
rect 649 -8 721 -4
rect 725 -8 744 -4
rect 748 -8 755 -4
rect 759 -8 858 -4
rect 862 -8 885 -4
rect 889 -8 931 -4
rect 935 -8 1000 -4
rect 1004 -8 1070 -4
rect 1074 -8 1140 -4
rect 1144 -8 1210 -4
rect 1214 -8 1293 -4
rect 1297 -8 1381 -4
rect 1385 -8 1514 -4
rect -42 -16 7 -12
rect 11 -16 79 -12
rect 83 -16 204 -12
rect 208 -16 352 -12
rect 356 -16 435 -12
rect 439 -16 509 -12
rect 513 -16 614 -12
rect 618 -16 686 -12
rect 690 -16 795 -12
rect 799 -16 823 -12
rect 827 -16 893 -12
rect 897 -16 939 -12
rect 943 -16 965 -12
rect 969 -16 1035 -12
rect 1039 -16 1105 -12
rect 1109 -16 1175 -12
rect 1179 -16 1258 -12
rect 1262 -16 1370 -12
rect 1374 -16 1514 -12
<< polycontact >>
rect -278 1785 -274 1789
rect -265 1775 -261 1779
rect -218 1774 -214 1778
rect -278 1767 -274 1771
rect -258 1751 -254 1755
rect -278 1739 -274 1743
rect 128 977 132 981
rect 150 997 154 1001
rect 1223 955 1227 959
rect 1287 853 1291 857
rect 1189 693 1193 697
rect 1287 603 1291 607
rect 1189 443 1193 447
rect 1287 353 1291 357
rect 1189 193 1193 197
rect 1287 103 1291 107
rect 1329 56 1333 60
<< m2contact >>
rect -265 1864 -261 1868
rect -313 1838 -309 1842
rect -277 1830 -273 1834
rect -258 1847 -254 1851
rect -218 1847 -214 1851
rect -204 1838 -200 1842
rect -173 1830 -169 1834
rect -155 1821 -151 1825
rect -111 1748 -107 1752
rect -103 1648 -99 1652
rect -110 875 -106 879
rect -95 1548 -91 1552
rect -102 750 -98 754
rect -87 1448 -83 1452
rect -94 625 -90 629
rect -79 1348 -75 1352
rect -86 500 -82 504
rect -71 1248 -67 1252
rect -78 375 -74 379
rect -63 1148 -59 1152
rect -70 250 -66 254
rect 1370 1675 1374 1679
rect 1287 1640 1291 1644
rect 1287 1619 1291 1623
rect 1370 1584 1374 1588
rect 1271 1573 1275 1577
rect 1287 1513 1291 1517
rect 1370 1470 1374 1474
rect 1287 1437 1291 1441
rect 1287 1416 1291 1420
rect 1370 1380 1374 1384
rect 1271 1370 1275 1374
rect 1287 1310 1291 1314
rect 1370 1266 1374 1270
rect 1287 1234 1291 1238
rect 1287 1213 1291 1217
rect 1370 1175 1374 1179
rect 1271 1167 1275 1171
rect -55 1048 -51 1052
rect -62 125 -58 129
rect 58 1012 62 1016
rect 98 1022 102 1026
rect 135 1012 139 1016
rect 192 1004 196 1008
rect 1287 1107 1291 1111
rect 1370 1061 1374 1065
rect 1287 1031 1291 1035
rect 1287 1010 1291 1014
rect 72 984 76 988
rect 1370 970 1374 974
rect 1271 964 1275 968
rect 1223 950 1227 954
rect 1287 904 1291 908
rect 1287 858 1291 862
rect 1370 841 1374 845
rect 1287 806 1291 810
rect 1287 785 1291 789
rect 1370 721 1374 725
rect 1271 714 1275 718
rect 1287 654 1291 658
rect 1287 608 1291 612
rect 1370 590 1374 594
rect 1287 556 1291 560
rect 1287 535 1291 539
rect 1370 471 1374 475
rect 1271 464 1275 468
rect 1287 404 1291 408
rect 1287 358 1291 362
rect 1370 340 1374 344
rect 1287 306 1291 310
rect 1287 285 1291 289
rect 1370 221 1374 225
rect 1271 214 1275 218
rect 1287 154 1291 158
rect 1287 108 1291 112
rect 1334 56 1338 60
rect 1287 35 1291 39
rect 1370 27 1374 31
rect -54 0 -50 4
rect 38 -8 42 -4
rect 121 -8 125 -4
rect 168 -8 172 -4
rect 317 -8 321 -4
rect 7 -16 11 -12
rect 79 -16 83 -12
rect 204 -16 208 -12
rect 393 -8 397 -4
rect 428 -8 432 -4
rect 352 -16 356 -12
rect 435 -16 439 -12
rect 509 -16 513 -12
rect 645 -8 649 -4
rect 721 -8 725 -4
rect 744 -8 748 -4
rect 755 -8 759 -4
rect 614 -16 618 -12
rect 686 -16 690 -12
rect 795 -16 799 -12
rect 858 -8 862 -4
rect 885 -8 889 -4
rect 931 -8 935 -4
rect 1000 -8 1004 -4
rect 1070 -8 1074 -4
rect 1140 -8 1144 -4
rect 1210 -8 1214 -4
rect 1293 -8 1297 -4
rect 1381 1596 1385 1600
rect 1381 1524 1385 1528
rect 1381 1391 1385 1395
rect 1381 1319 1385 1323
rect 1381 1186 1385 1190
rect 1381 1114 1385 1118
rect 1381 981 1385 985
rect 1381 909 1385 913
rect 1381 761 1385 765
rect 1381 689 1385 693
rect 1381 511 1385 515
rect 1381 439 1385 443
rect 1381 261 1385 265
rect 1381 189 1385 193
rect 1381 87 1385 91
rect 1381 -8 1385 -4
rect 823 -16 827 -12
rect 893 -16 897 -12
rect 939 -16 943 -12
rect 965 -16 969 -12
rect 1035 -16 1039 -12
rect 1105 -16 1109 -12
rect 1175 -16 1179 -12
rect 1258 -16 1262 -12
rect 1370 -16 1374 -12
use ir_register  InstructionRegister
timestamp 1434186535
transform 1 0 -218 0 1 957
box 0 0 103 848
use additiveAccumulatorController  additiveAccumulatorController_0
timestamp 1434090485
transform 1 0 151 0 1 1222
box -91 -192 83 -98
use input_register  input_register_0
timestamp 1434158754
transform 1 0 0 0 1 0
box -42 0 48 1028
use adder  reg_a
timestamp 1434092755
transform 1 0 51 0 1 0
box 0 0 270 1026
use fblock  reg_l
timestamp 1434148540
transform 1 0 324 0 1 0
box 0 0 232 1120
use shifter  reg_s
timestamp 1434151676
transform 1 0 557 0 1 0
box -4 0 111 1064
use pwm  reg_p
timestamp 1434158785
transform 1 0 671 0 1 0
box 0 0 276 1091
use register  reg4
timestamp 1434142685
transform 1 0 950 0 1 0
box 0 0 67 1032
use register  reg5
timestamp 1434142685
transform 1 0 1020 0 1 0
box 0 0 67 1032
use register  reg6
timestamp 1434142685
transform 1 0 1090 0 1 0
box 0 0 67 1032
use register  reg7
timestamp 1434142685
transform 1 0 1160 0 1 0
box 0 0 67 1032
use pcregister  pcregister_0
timestamp 1434174971
transform 1 0 1237 0 1 0
box -38 0 140 1823
use pcIncrementor  pcIncrementor_0
timestamp 1434180000
transform -1 0 1812 0 1 0
box 298 0 422 1679
<< labels >>
rlabel metal2 -216 1832 -216 1832 3 Vdd
rlabel metal2 -215 1840 -215 1840 4 GND
rlabel metal2 -311 1849 -311 1849 1 phi0
rlabel metal2 -311 1858 -311 1858 1 phi0_
rlabel metal2 -311 1866 -311 1866 1 phi1
rlabel metal2 -311 1874 -311 1874 5 phi1_
rlabel metal2 -311 1882 -311 1882 5 RESET
rlabel metal2 -303 1822 -303 1822 1 RESET_
<< end >>
