magic
tech scmos
timestamp 1434160103
<< polysilicon >>
rect -16 23 -14 25
rect 18 23 28 25
rect -16 19 -14 21
rect 18 19 24 21
rect 22 13 24 19
rect 1 11 24 13
rect 1 7 3 11
rect 26 8 28 23
rect -7 5 3 7
rect 1 1 3 5
rect 18 6 28 8
rect 18 4 19 6
rect 17 1 19 4
rect 1 -9 3 -7
rect 17 -9 19 -7
<< ndiffusion >>
rect 0 -7 1 1
rect 3 -7 4 1
rect 16 -7 17 1
rect 19 -7 20 1
<< pdiffusion >>
rect -14 25 18 26
rect -14 21 18 23
rect -14 18 18 19
<< metal1 >>
rect 18 14 24 18
rect -4 1 -1 14
rect 21 8 24 14
rect 8 4 14 7
rect 21 5 38 8
rect 8 1 12 4
rect 21 1 24 5
<< ntransistor >>
rect 1 -7 3 1
rect 17 -7 19 1
<< ptransistor >>
rect -14 23 18 25
rect -14 19 18 21
<< polycontact >>
rect -11 5 -7 9
rect 14 4 18 8
<< ndcontact >>
rect -4 -7 0 1
rect 4 -7 8 1
rect 12 -7 16 1
rect 20 -7 24 1
<< pdcontact >>
rect -14 26 18 30
rect -14 14 18 18
<< psubstratepcontact >>
rect 8 -7 12 1
<< nsubstratencontact >>
rect -14 30 18 34
<< labels >>
rlabel polycontact -9 7 -9 7 3 cin
rlabel metal1 36 6 36 6 7 cout
<< end >>
