magic
tech scmos
timestamp 1434159111
<< polysilicon >>
rect -14 5 -12 7
rect 4 5 8 7
rect 6 -15 8 5
rect -8 -17 -6 -15
rect 2 -17 8 -15
<< ndiffusion >>
rect -6 -15 2 -14
rect -6 -18 2 -17
<< pdiffusion >>
rect -12 7 4 8
rect -12 4 4 5
<< metal1 >>
rect -2 -10 2 0
<< ntransistor >>
rect -6 -17 2 -15
<< ptransistor >>
rect -12 5 4 7
<< ndcontact >>
rect -6 -14 2 -10
rect -6 -22 2 -18
<< pdcontact >>
rect -12 8 4 12
rect -12 0 4 4
<< psubstratepcontact >>
rect -6 -26 2 -22
<< nsubstratencontact >>
rect -12 12 4 16
<< end >>
