magic
tech scmos
timestamp 1434144344
<< polysilicon >>
rect -13 38 37 40
rect -13 24 -11 38
rect 3 33 14 35
rect 3 32 5 33
rect -9 30 -7 32
rect 1 30 5 32
rect -16 22 -7 24
rect 1 22 3 24
rect 12 21 14 33
rect 16 30 27 32
rect 31 30 33 32
rect 16 17 18 30
rect 35 24 37 38
rect 25 22 27 24
rect 31 22 37 24
rect 16 8 18 13
rect -16 6 -7 8
rect 1 6 18 8
rect 25 6 27 8
rect 31 6 40 8
rect 19 3 27 4
rect -9 -2 -7 0
rect 1 -2 7 0
rect 17 2 27 3
rect 31 2 33 4
rect 17 1 21 2
rect 5 -5 7 -2
rect 35 -5 37 6
rect 5 -7 37 -5
<< ndiffusion >>
rect 27 32 31 33
rect 27 29 31 30
rect 27 24 31 25
rect 27 21 31 22
rect 15 13 16 17
rect 18 13 19 17
rect 27 8 31 9
rect 27 4 31 6
rect 27 1 31 2
<< pdiffusion >>
rect -7 32 1 33
rect -7 29 1 30
rect -7 24 1 25
rect -7 21 1 22
rect -7 8 1 9
rect -7 5 1 6
rect -7 0 1 1
rect -7 -3 1 -2
<< metal1 >>
rect 11 37 14 43
rect -13 33 -7 36
rect 1 34 27 37
rect 31 34 37 37
rect -13 -4 -10 33
rect 4 30 6 31
rect 1 27 6 30
rect 10 30 16 31
rect 10 29 18 30
rect 10 28 27 29
rect 13 27 27 28
rect 1 26 4 27
rect 15 26 27 27
rect 12 20 14 23
rect 11 17 14 20
rect 1 13 2 17
rect 23 13 27 17
rect 11 4 14 13
rect 1 3 17 4
rect 1 1 13 3
rect -13 -7 -7 -4
rect 20 -8 23 13
rect 34 0 37 34
rect 40 10 43 26
rect 31 -3 37 0
rect 20 -11 43 -8
<< metal2 >>
rect 10 29 18 30
rect 10 26 40 29
rect -16 13 2 17
<< ntransistor >>
rect 27 30 31 32
rect 27 22 31 24
rect 16 13 18 17
rect 27 6 31 8
rect 27 2 31 4
<< ptransistor >>
rect -7 30 1 32
rect -7 22 1 24
rect -7 6 1 8
rect -7 -2 1 0
<< polycontact >>
rect -20 22 -16 26
rect 8 20 12 24
rect -20 4 -16 8
rect 40 6 44 10
rect 13 -1 17 3
<< ndcontact >>
rect 27 33 31 37
rect 27 25 31 29
rect 27 17 31 21
rect 11 13 15 17
rect 19 13 23 17
rect 27 9 31 13
rect 27 -3 31 1
<< pdcontact >>
rect -7 33 1 37
rect -7 25 1 29
rect -7 17 1 21
rect -7 9 1 13
rect -7 1 1 5
rect -7 -7 1 -3
<< m2contact >>
rect -20 13 -16 17
rect 6 27 10 31
rect 2 13 6 17
rect 40 26 44 30
<< psubstratepcontact >>
rect 27 13 31 17
<< nsubstratencontact >>
rect -7 13 1 17
<< labels >>
rlabel polysilicon -8 23 -8 23 3 b
rlabel polysilicon -8 31 -8 31 3 a_
rlabel polysilicon -8 7 -8 7 3 a
rlabel polysilicon -8 -1 -8 -1 3 b_
rlabel polysilicon 26 3 26 3 1 a_
rlabel metal1 12 42 12 42 5 xor
rlabel metal1 41 -10 41 -10 8 GND
rlabel m2contact -18 15 -18 15 3 Vdd
rlabel polycontact -18 6 -18 6 3 a
rlabel polycontact -18 24 -18 24 3 b
<< end >>
