magic
tech scmos
timestamp 1432009782
<< metal1 >>
rect 307 1270 438 1274
rect 280 1262 288 1266
rect 140 1258 288 1262
rect 67 909 71 1252
rect 140 1218 143 1258
rect 292 1254 295 1266
rect 300 1263 303 1266
rect 179 1250 295 1254
rect 89 1120 93 1187
rect 179 1152 183 1250
rect 307 1246 311 1270
rect 435 1263 438 1266
rect 443 1257 446 1272
rect 273 1242 311 1246
rect 315 1253 446 1257
rect 187 1199 191 1222
rect 179 1103 183 1107
rect 273 1067 277 1242
rect 315 1238 319 1253
rect 282 1234 319 1238
rect 282 1035 286 1234
rect 450 1230 458 1274
rect 309 1226 458 1230
rect 290 997 293 1063
rect 164 992 167 995
rect 171 992 174 995
rect 297 988 301 1040
rect 309 1026 313 1226
rect 320 1218 549 1222
rect 320 1044 324 1218
rect 554 1214 558 1251
rect 329 1210 558 1214
rect 329 1081 333 1210
rect 570 1206 574 1251
rect 337 1202 574 1206
rect 337 1180 341 1202
rect 578 1198 582 1251
rect 390 1022 394 1195
rect 553 1194 582 1198
rect 279 984 301 988
rect 553 987 556 1194
rect 586 1190 590 1251
rect 560 1186 590 1190
rect 560 1084 564 1186
rect 594 1183 598 1251
rect 572 1179 598 1183
rect 602 1095 606 1251
rect 610 1191 614 1251
rect 651 1042 695 1046
rect 651 1032 655 1042
rect 691 909 695 1042
<< metal2 >>
rect 103 1266 106 1269
rect 119 1266 122 1269
rect 135 1266 138 1269
rect 151 1266 154 1269
rect 167 1256 170 1269
rect 71 1252 170 1256
rect 183 1226 186 1269
rect 263 1266 485 1270
rect 199 1234 202 1266
rect 215 1243 218 1266
rect 231 1252 234 1266
rect 247 1262 250 1266
rect 490 1262 493 1267
rect 247 1258 493 1262
rect 498 1252 501 1267
rect 231 1248 501 1252
rect 506 1243 509 1266
rect 215 1239 509 1243
rect 514 1234 517 1266
rect 522 1263 525 1266
rect 530 1263 533 1266
rect 538 1263 541 1266
rect 199 1230 517 1234
rect 546 1226 549 1266
rect 554 1255 557 1266
rect 570 1255 573 1266
rect 578 1255 581 1266
rect 586 1255 589 1266
rect 594 1255 597 1266
rect 602 1255 605 1266
rect 610 1255 613 1266
rect 183 1222 187 1226
rect 618 1218 621 1266
rect 121 1214 621 1218
rect 191 1195 390 1199
rect 93 1187 610 1191
rect 208 1176 337 1180
rect 481 1179 568 1183
rect 93 1116 125 1120
rect 23 1091 602 1095
rect 23 1060 27 1091
rect 208 1077 329 1081
rect 481 1080 560 1084
rect 277 1063 290 1067
rect 301 1040 320 1044
rect 0 964 4 968
rect 247 933 251 937
rect 71 905 691 909
rect 0 839 4 843
rect 247 808 251 812
rect 0 714 4 718
rect 247 683 251 687
rect 0 589 4 593
rect 247 558 251 562
rect 0 464 4 468
rect 247 433 251 437
rect 0 339 4 343
rect 247 308 251 312
rect 0 214 4 218
rect 247 183 251 187
rect 0 89 4 93
rect 247 58 251 62
rect 11 8 15 12
rect 11 0 15 4
<< m2contact >>
rect 67 1252 71 1256
rect 24 964 28 968
rect 89 1187 93 1191
rect 187 1222 191 1226
rect 187 1195 191 1199
rect 179 1148 183 1152
rect 89 1116 93 1120
rect 273 1063 277 1067
rect 554 1251 558 1255
rect 282 1031 286 1035
rect 290 1063 294 1067
rect 289 993 293 997
rect 297 1040 301 1044
rect 545 1222 549 1226
rect 570 1251 574 1255
rect 578 1251 582 1255
rect 337 1176 341 1180
rect 390 1195 394 1199
rect 329 1077 333 1081
rect 320 1040 324 1044
rect 586 1251 590 1255
rect 594 1251 598 1255
rect 568 1179 572 1183
rect 602 1251 606 1255
rect 610 1251 614 1255
rect 610 1187 614 1191
rect 602 1091 606 1095
rect 560 1080 564 1084
rect 67 905 71 909
rect 691 905 695 909
rect 24 839 28 843
rect 24 714 28 718
rect 24 589 28 593
rect 24 464 28 468
rect 24 339 28 343
rect 24 214 28 218
rect 24 89 28 93
use divide_ctl  divide_ctl_0
timestamp 1432009782
transform 1 0 64 0 1 1843
box 0 -577 579 30
use divide_datapath  divide_datapath_0
timestamp 1431680467
transform 1 0 433 0 1 0
box -433 0 259 1218
<< labels >>
rlabel metal2 11 0 15 4 1 Vdd
rlabel metal2 11 8 15 12 1 GND
rlabel metal2 0 89 4 93 3 dout0
rlabel m2contact 24 89 28 93 1 din0
rlabel metal2 0 214 4 218 3 dout1
rlabel m2contact 24 214 28 218 1 din1
rlabel metal2 0 339 4 343 3 dout2
rlabel m2contact 24 339 28 343 1 din2
rlabel metal2 0 464 4 468 3 dout3
rlabel m2contact 24 464 28 468 1 din3
rlabel metal2 0 589 4 593 3 dout4
rlabel m2contact 24 589 28 593 1 din4
rlabel metal2 0 714 4 718 3 dout5
rlabel m2contact 24 714 28 718 1 din5
rlabel metal2 0 839 4 843 3 dout6
rlabel m2contact 24 839 28 843 1 din6
rlabel metal2 0 964 4 968 3 dout7
rlabel m2contact 24 964 28 968 1 din7
rlabel metal2 103 1266 106 1269 1 RESET
rlabel metal2 119 1266 122 1269 1 req_d
rlabel metal2 135 1266 138 1269 1 req_v
rlabel metal2 151 1266 154 1269 1 ack_out
rlabel metal1 292 1263 295 1266 1 phi0
rlabel metal1 300 1263 303 1266 1 phi0_
rlabel metal1 435 1263 438 1266 1 phi1_
rlabel metal1 443 1263 446 1266 1 phi1
rlabel metal2 522 1263 525 1266 1 ack_in
rlabel metal2 530 1263 533 1266 1 req_Q
rlabel metal2 538 1263 541 1266 1 req_R
rlabel metal2 167 1252 170 1256 1 icarry
rlabel metal2 183 1254 186 1258 1 scarry
rlabel metal2 247 933 251 937 1 acc7
rlabel metal2 247 808 251 812 1 acc6
rlabel metal2 247 683 251 687 1 acc5
rlabel metal2 247 558 251 562 1 acc4
rlabel metal2 247 433 251 437 1 acc3
rlabel metal2 247 308 251 312 1 acc2
rlabel metal2 247 183 251 187 1 acc1
rlabel metal2 247 58 251 62 1 acc0
rlabel metal1 171 992 174 995 1 accw
rlabel metal1 164 992 167 995 1 accw_
<< end >>
