magic
tech scmos
timestamp 1433955363
<< polysilicon >>
rect -40 14 -19 16
rect 7 14 26 16
rect 5 2 7 4
rect -33 -2 -19 0
rect 7 -2 19 0
rect 7 -46 9 -38
rect -26 -60 -3 -58
rect 5 -60 7 -58
<< pdiffusion >>
rect -3 -58 5 -57
rect -3 -61 5 -60
<< metal1 >>
rect -44 17 -41 21
rect -44 -65 -41 13
rect -37 1 -34 21
rect -37 -65 -34 -3
rect -30 -57 -27 21
rect -23 9 -20 21
rect -9 18 -7 21
rect -23 5 -17 9
rect 13 9 16 21
rect -23 -31 -20 5
rect -10 -20 -6 7
rect 5 5 16 9
rect 6 -21 9 -18
rect 13 -31 16 5
rect 20 1 23 21
rect 27 17 30 21
rect -23 -35 -17 -31
rect 11 -35 16 -31
rect -30 -65 -27 -61
rect -23 -65 -20 -35
rect -10 -43 -6 -39
rect 2 -50 6 -47
rect 2 -53 5 -50
rect 13 -61 16 -35
rect 5 -65 16 -61
rect 20 -65 23 -3
rect 27 -65 30 13
<< ptransistor >>
rect -3 -60 5 -58
<< polycontact >>
rect -44 13 -40 17
rect 26 13 30 17
rect -10 7 -6 11
rect -37 -3 -33 1
rect 19 -3 23 1
rect 6 -50 10 -46
rect -30 -61 -26 -57
<< pdcontact >>
rect -3 -57 5 -53
rect -3 -65 5 -61
use latch  latch_1
timestamp 1430426212
transform 0 1 -17 1 0 11
box -6 -2 10 24
use latch  latch_0
timestamp 1430426212
transform 0 1 -17 -1 0 3
box -6 -2 10 24
use staticizer  staticizer_0
timestamp 1430428783
transform 0 1 -21 -1 0 -31
box -19 2 12 32
<< labels >>
rlabel metal1 -10 -43 -6 -39 1 cnt
rlabel metal1 -9 18 -7 21 5 out
rlabel polysilicon 5 2 7 4 7 in
rlabel metal1 -23 18 -20 21 5 GND
rlabel metal1 13 18 16 21 5 Vdd
rlabel metal1 20 18 23 21 5 w_
rlabel metal1 -30 18 -27 21 5 reset
rlabel metal1 -37 18 -34 21 5 w
rlabel metal1 -44 18 -41 21 4 r
rlabel metal1 27 18 30 21 6 r_
rlabel metal1 6 -21 9 -18 1 cnt_
<< end >>
