magic
tech scmos
timestamp 1434175533
<< polysilicon >>
rect -48 23 -46 25
rect 18 23 28 25
rect -48 19 -46 21
rect 18 19 24 21
rect 22 13 24 19
rect 1 11 24 13
rect 1 7 3 11
rect 26 8 28 23
rect -7 5 3 7
rect 1 1 3 5
rect 17 6 28 8
rect 17 1 19 6
rect 1 -17 3 -15
rect 17 -17 19 -15
<< ndiffusion >>
rect 0 -15 1 1
rect 3 -15 4 1
rect 16 -15 17 1
rect 19 -15 20 1
<< pdiffusion >>
rect -46 25 18 26
rect -46 21 18 23
rect -46 18 18 19
<< metal1 >>
rect 18 14 24 18
rect -76 5 -11 9
rect -4 1 -1 14
rect 21 8 24 14
rect 21 5 35 8
rect 21 1 24 5
<< ntransistor >>
rect 1 -15 3 1
rect 17 -15 19 1
<< ptransistor >>
rect -46 23 18 25
rect -46 19 18 21
<< polycontact >>
rect -11 5 -7 9
<< ndcontact >>
rect -4 -15 0 1
rect 4 -15 8 1
rect 12 -15 16 1
rect 20 -15 24 1
<< pdcontact >>
rect -46 26 18 30
rect -46 14 18 18
<< psubstratepcontact >>
rect 8 -15 12 1
<< nsubstratencontact >>
rect -46 30 18 34
<< labels >>
rlabel polycontact -9 7 -9 7 3 cin
<< end >>
